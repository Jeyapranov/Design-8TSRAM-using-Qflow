magic
tech scmos
timestamp 1751994658
<< metal1 >>
rect 888 1703 890 1707
rect 894 1703 897 1707
rect 901 1703 904 1707
rect 1062 1678 1074 1681
rect 1070 1677 1074 1678
rect 406 1668 414 1671
rect 1038 1668 1046 1671
rect 6 1658 33 1661
rect 198 1658 206 1661
rect 406 1658 425 1661
rect 878 1658 886 1661
rect 1038 1658 1057 1661
rect 1122 1658 1129 1661
rect 1366 1652 1369 1662
rect 1519 1658 1537 1661
rect 1746 1658 1753 1661
rect 675 1638 678 1642
rect 368 1603 370 1607
rect 374 1603 377 1607
rect 381 1603 384 1607
rect 1384 1603 1386 1607
rect 1390 1603 1393 1607
rect 1397 1603 1400 1607
rect 210 1588 211 1592
rect 930 1588 931 1592
rect 1790 1588 1798 1591
rect 538 1578 539 1582
rect 94 1568 102 1571
rect 1013 1568 1014 1572
rect 1154 1568 1157 1572
rect 110 1548 129 1551
rect 222 1548 241 1551
rect 550 1548 569 1551
rect 638 1548 657 1551
rect 790 1542 793 1551
rect 942 1548 961 1551
rect 982 1548 1001 1551
rect 1238 1548 1257 1551
rect 1326 1548 1345 1551
rect 122 1538 129 1541
rect 246 1538 254 1541
rect 362 1538 370 1541
rect 578 1538 585 1541
rect 638 1538 646 1541
rect 1326 1538 1334 1541
rect 246 1528 249 1538
rect 454 1531 458 1533
rect 454 1528 465 1531
rect 470 1528 489 1531
rect 574 1528 577 1538
rect 670 1531 674 1533
rect 662 1528 674 1531
rect 686 1532 690 1536
rect 594 1518 595 1522
rect 888 1503 890 1507
rect 894 1503 897 1507
rect 901 1503 904 1507
rect 682 1488 689 1491
rect 1018 1488 1019 1492
rect 1382 1488 1393 1491
rect 110 1478 129 1481
rect 204 1478 206 1482
rect 270 1478 282 1481
rect 414 1478 433 1481
rect 862 1478 890 1481
rect 1382 1481 1385 1488
rect 1206 1478 1218 1481
rect 1366 1478 1385 1481
rect 278 1477 282 1478
rect 886 1477 890 1478
rect 1214 1477 1218 1478
rect 246 1468 254 1471
rect 660 1468 670 1471
rect 838 1468 846 1471
rect 1030 1468 1046 1471
rect 1302 1468 1310 1471
rect 1510 1471 1513 1481
rect 1590 1478 1609 1481
rect 1510 1468 1529 1471
rect 126 1458 129 1468
rect 166 1458 186 1461
rect 246 1458 265 1461
rect 838 1458 857 1461
rect 1038 1458 1046 1461
rect 1078 1458 1086 1461
rect 1094 1458 1113 1461
rect 1182 1458 1201 1461
rect 1358 1458 1366 1461
rect 1534 1458 1542 1461
rect 182 1456 186 1458
rect 590 1448 609 1451
rect 186 1438 201 1441
rect 574 1438 590 1441
rect 368 1403 370 1407
rect 374 1403 377 1407
rect 381 1403 384 1407
rect 1384 1403 1386 1407
rect 1390 1403 1393 1407
rect 1397 1403 1400 1407
rect 1746 1388 1747 1392
rect 266 1368 281 1371
rect 258 1358 265 1361
rect 342 1358 353 1361
rect 710 1358 721 1361
rect 1642 1358 1649 1361
rect 718 1352 721 1358
rect 230 1348 249 1351
rect 430 1348 438 1351
rect 882 1348 913 1351
rect 310 1341 313 1348
rect 1094 1348 1102 1351
rect 1110 1348 1129 1351
rect 1266 1348 1273 1351
rect 1282 1348 1289 1351
rect 1330 1348 1337 1351
rect 1366 1348 1374 1351
rect 1502 1348 1545 1351
rect 1634 1348 1657 1351
rect 1782 1351 1785 1358
rect 1762 1348 1777 1351
rect 1782 1348 1793 1351
rect 302 1338 313 1341
rect 502 1338 521 1341
rect 882 1338 905 1341
rect 1282 1338 1289 1341
rect 372 1328 382 1331
rect 518 1328 521 1338
rect 1254 1331 1258 1333
rect 1254 1328 1265 1331
rect 1782 1328 1785 1338
rect 650 1318 651 1322
rect 669 1318 670 1322
rect 805 1318 806 1322
rect 857 1318 886 1321
rect 1698 1318 1699 1322
rect 888 1303 890 1307
rect 894 1303 897 1307
rect 901 1303 904 1307
rect 29 1288 30 1292
rect 793 1288 798 1292
rect 394 1278 395 1282
rect 458 1278 459 1282
rect 762 1278 769 1281
rect 910 1278 937 1281
rect 1046 1278 1065 1281
rect 1306 1278 1307 1282
rect 1382 1278 1390 1281
rect 1486 1278 1494 1281
rect 910 1277 914 1278
rect 1206 1272 1209 1278
rect 102 1268 110 1271
rect 130 1268 138 1271
rect 770 1268 777 1271
rect 954 1268 961 1271
rect 1206 1268 1210 1272
rect 1274 1268 1281 1271
rect 1370 1268 1377 1271
rect 1410 1268 1417 1271
rect 1478 1268 1486 1271
rect 54 1258 62 1261
rect 102 1258 121 1261
rect 406 1258 425 1261
rect 470 1258 489 1261
rect 854 1258 862 1261
rect 942 1258 961 1261
rect 998 1261 1001 1268
rect 998 1258 1009 1261
rect 1554 1258 1561 1261
rect 1634 1258 1641 1261
rect 206 1252 210 1257
rect 694 1241 697 1251
rect 678 1238 697 1241
rect 910 1238 934 1241
rect 678 1228 681 1238
rect 368 1203 370 1207
rect 374 1203 377 1207
rect 381 1203 384 1207
rect 1384 1203 1386 1207
rect 1390 1203 1393 1207
rect 1397 1203 1400 1207
rect 29 1168 30 1172
rect 1374 1168 1390 1171
rect 818 1158 825 1161
rect 550 1153 554 1158
rect 54 1148 62 1151
rect 274 1148 281 1151
rect 446 1148 465 1151
rect 678 1148 697 1151
rect 886 1148 921 1151
rect 930 1148 937 1151
rect 1102 1148 1121 1151
rect 1358 1148 1377 1151
rect 1646 1148 1665 1151
rect 1738 1148 1761 1151
rect 370 1138 393 1141
rect 738 1138 753 1141
rect 886 1138 910 1141
rect 938 1138 945 1141
rect 1358 1138 1366 1141
rect 1674 1138 1681 1141
rect 1726 1138 1753 1141
rect 830 1132 833 1138
rect 190 1128 209 1131
rect 342 1128 361 1131
rect 830 1128 838 1132
rect 1382 1128 1401 1131
rect 1634 1128 1635 1132
rect 1670 1128 1673 1138
rect 709 1118 710 1122
rect 769 1118 790 1121
rect 1398 1121 1401 1128
rect 1398 1118 1409 1121
rect 1690 1118 1691 1122
rect 888 1103 890 1107
rect 894 1103 897 1107
rect 901 1103 904 1107
rect 502 1088 510 1091
rect 1390 1088 1401 1091
rect 126 1078 145 1081
rect 218 1078 234 1081
rect 230 1074 234 1078
rect 590 1071 593 1081
rect 1398 1081 1401 1088
rect 1398 1078 1417 1081
rect 1702 1078 1714 1081
rect 574 1068 593 1071
rect 822 1071 825 1078
rect 1710 1077 1714 1078
rect 786 1068 793 1071
rect 812 1068 825 1071
rect 834 1068 849 1071
rect 894 1068 910 1071
rect 1198 1068 1210 1071
rect 1422 1068 1433 1071
rect 246 1058 257 1061
rect 402 1058 409 1061
rect 438 1058 457 1061
rect 654 1061 657 1068
rect 654 1058 665 1061
rect 722 1058 737 1061
rect 826 1058 841 1061
rect 1050 1058 1057 1061
rect 1086 1058 1094 1061
rect 1430 1062 1433 1068
rect 1334 1058 1342 1061
rect 1482 1058 1489 1061
rect 1694 1058 1702 1061
rect 246 1057 250 1058
rect 474 1048 481 1051
rect 698 1038 701 1042
rect 1730 1038 1733 1042
rect 368 1003 370 1007
rect 374 1003 377 1007
rect 381 1003 384 1007
rect 1384 1003 1386 1007
rect 1390 1003 1393 1007
rect 1397 1003 1400 1007
rect 1125 988 1126 992
rect 770 968 773 972
rect 110 948 129 951
rect 306 948 321 951
rect 558 948 574 951
rect 694 948 713 951
rect 914 948 921 951
rect 1050 948 1065 951
rect 1106 948 1113 951
rect 1638 948 1646 951
rect 122 938 129 941
rect 190 938 206 941
rect 214 938 233 941
rect 706 938 713 941
rect 94 931 98 933
rect 94 928 105 931
rect 230 928 233 938
rect 678 931 682 933
rect 678 928 689 931
rect 1154 928 1161 931
rect 1166 928 1182 931
rect 1654 931 1658 933
rect 1646 928 1658 931
rect 189 918 190 922
rect 370 918 377 921
rect 858 918 865 921
rect 888 903 890 907
rect 894 903 897 907
rect 901 903 904 907
rect 246 888 257 891
rect 458 888 459 892
rect 650 888 652 892
rect 909 888 910 892
rect 1205 888 1206 892
rect 254 882 257 888
rect 138 878 145 881
rect 150 871 153 878
rect 122 868 137 871
rect 150 868 161 871
rect 286 868 294 871
rect 102 858 105 868
rect 134 858 137 868
rect 174 861 177 868
rect 166 858 177 861
rect 310 861 313 871
rect 394 868 417 871
rect 590 871 593 881
rect 690 878 697 882
rect 710 878 729 881
rect 942 878 961 881
rect 1013 878 1014 882
rect 1126 878 1137 881
rect 1366 878 1385 881
rect 1390 878 1406 881
rect 1614 878 1633 881
rect 694 872 697 878
rect 1126 877 1130 878
rect 1638 872 1641 881
rect 590 868 609 871
rect 802 868 817 871
rect 974 868 990 871
rect 1710 868 1737 871
rect 290 858 313 861
rect 346 856 361 859
rect 670 858 681 861
rect 862 858 897 861
rect 926 858 934 861
rect 1714 858 1745 861
rect 670 856 674 858
rect 678 852 681 858
rect 342 848 350 851
rect 1230 848 1238 851
rect 370 838 377 841
rect 382 818 390 821
rect 368 803 370 807
rect 374 803 377 807
rect 381 803 384 807
rect 1384 803 1386 807
rect 1390 803 1393 807
rect 1397 803 1400 807
rect 222 768 230 771
rect 578 768 585 771
rect 750 768 766 771
rect 770 768 777 771
rect 222 766 226 768
rect 766 752 770 754
rect 150 748 169 751
rect 366 748 401 751
rect 634 748 641 751
rect 686 748 705 751
rect 914 748 921 751
rect 1290 748 1305 751
rect 1362 748 1374 751
rect 1686 748 1694 751
rect 110 738 121 741
rect 162 738 169 741
rect 378 738 401 741
rect 798 738 814 741
rect 986 738 993 741
rect 998 738 1006 741
rect 1146 738 1158 741
rect 1286 738 1294 741
rect 110 732 113 738
rect 350 731 354 733
rect 350 728 361 731
rect 798 728 801 738
rect 1022 728 1030 731
rect 1038 728 1046 731
rect 1142 728 1158 731
rect 888 703 890 707
rect 894 703 897 707
rect 901 703 904 707
rect 874 688 875 692
rect 914 688 921 691
rect 222 668 238 671
rect 262 668 270 671
rect 366 668 382 671
rect 490 668 497 671
rect 510 671 513 681
rect 602 678 609 681
rect 614 678 633 681
rect 790 678 801 681
rect 1334 678 1345 681
rect 1674 678 1681 681
rect 790 677 794 678
rect 1334 677 1338 678
rect 510 668 529 671
rect 546 668 561 671
rect 818 668 825 671
rect 866 668 873 671
rect 886 668 910 671
rect 1034 668 1041 671
rect 1506 668 1518 671
rect 1546 668 1553 671
rect 78 658 86 661
rect 310 658 318 661
rect 654 658 662 661
rect 806 658 825 661
rect 1022 658 1041 661
rect 1230 658 1238 661
rect 1346 658 1353 661
rect 1566 658 1582 661
rect 1586 658 1593 661
rect 1738 658 1753 661
rect 598 651 601 658
rect 590 648 601 651
rect 1434 648 1438 652
rect 1370 618 1371 622
rect 1642 618 1643 622
rect 368 603 370 607
rect 374 603 377 607
rect 381 603 384 607
rect 1384 603 1386 607
rect 1390 603 1393 607
rect 1397 603 1400 607
rect 717 588 718 592
rect 234 568 241 571
rect 398 568 406 571
rect 1374 558 1382 561
rect 1628 557 1630 561
rect 54 548 62 551
rect 410 548 425 551
rect 494 548 505 551
rect 706 548 713 551
rect 766 548 785 551
rect 794 548 801 551
rect 494 542 497 548
rect 1110 548 1129 551
rect 1734 548 1742 551
rect 62 538 78 541
rect 226 538 233 541
rect 510 538 518 541
rect 690 538 697 541
rect 790 538 798 541
rect 802 538 809 541
rect 974 538 993 541
rect 1122 538 1129 541
rect 1386 538 1409 541
rect 62 528 65 538
rect 278 528 297 531
rect 790 528 793 538
rect 974 528 977 538
rect 1254 528 1262 531
rect 29 518 30 522
rect 754 518 755 522
rect 888 503 890 507
rect 894 503 897 507
rect 901 503 904 507
rect 194 488 195 492
rect 894 488 902 491
rect 1005 488 1006 492
rect 334 478 350 481
rect 654 478 665 481
rect 938 478 939 482
rect 1390 478 1406 481
rect 178 468 185 471
rect 310 468 318 471
rect 570 468 582 471
rect 590 468 606 471
rect 662 471 665 478
rect 662 468 670 471
rect 686 468 697 471
rect 766 468 769 478
rect 1018 468 1033 471
rect 1274 468 1281 471
rect 310 458 329 461
rect 686 462 689 468
rect 642 458 662 461
rect 742 458 750 461
rect 950 458 969 461
rect 1230 458 1246 461
rect 1370 458 1385 461
rect 1618 458 1625 461
rect 686 448 697 451
rect 875 438 878 442
rect 368 403 370 407
rect 374 403 377 407
rect 381 403 384 407
rect 1384 403 1386 407
rect 1390 403 1393 407
rect 1397 403 1400 407
rect 813 388 814 392
rect 1210 388 1211 392
rect 1461 388 1462 392
rect 1770 388 1771 392
rect 470 371 473 381
rect 454 368 473 371
rect 454 358 457 368
rect 646 361 649 368
rect 638 358 649 361
rect 1434 358 1449 361
rect 494 352 498 354
rect 318 348 337 351
rect 382 348 417 351
rect 582 348 590 351
rect 730 348 745 351
rect 766 348 777 351
rect 862 348 870 351
rect 918 348 937 351
rect 774 342 777 348
rect 1146 348 1161 351
rect 1598 348 1617 351
rect 1686 348 1694 351
rect 106 338 113 341
rect 614 338 622 341
rect 306 328 307 332
rect 626 328 633 331
rect 778 328 785 331
rect 1054 328 1073 331
rect 1566 331 1570 333
rect 1566 328 1577 331
rect 888 303 890 307
rect 894 303 897 307
rect 901 303 904 307
rect 189 288 190 292
rect 532 288 534 292
rect 653 288 654 292
rect 1165 288 1166 292
rect 1253 288 1254 292
rect 1421 288 1422 292
rect 94 278 105 281
rect 922 278 937 281
rect 1058 278 1066 281
rect 94 277 98 278
rect 1062 277 1066 278
rect 122 268 129 271
rect 378 268 393 271
rect 418 268 425 271
rect 438 268 446 271
rect 110 258 129 261
rect 410 258 417 261
rect 550 261 553 271
rect 626 268 633 271
rect 662 268 673 271
rect 762 268 785 271
rect 798 268 809 271
rect 954 268 961 271
rect 1030 268 1038 271
rect 1214 268 1222 271
rect 1270 271 1274 274
rect 1266 268 1274 271
rect 1438 271 1441 278
rect 1430 268 1441 271
rect 1746 268 1753 271
rect 798 262 801 268
rect 550 258 569 261
rect 606 258 625 261
rect 754 258 774 261
rect 942 258 961 261
rect 990 258 998 261
rect 1030 258 1049 261
rect 1214 258 1233 261
rect 1382 258 1406 261
rect 1486 258 1494 261
rect 1638 258 1646 261
rect 1774 258 1793 261
rect 406 248 409 258
rect 574 248 585 251
rect 798 248 809 251
rect 1774 248 1777 258
rect 498 238 529 241
rect 602 238 609 241
rect 368 203 370 207
rect 374 203 377 207
rect 381 203 384 207
rect 1384 203 1386 207
rect 1390 203 1393 207
rect 1397 203 1400 207
rect 1461 188 1462 192
rect 1650 188 1651 192
rect 146 168 149 172
rect 54 158 62 161
rect 1138 158 1145 161
rect 1702 158 1710 161
rect 1722 158 1729 161
rect 254 148 273 151
rect 338 148 345 151
rect 430 148 457 151
rect 622 148 641 151
rect 918 148 937 151
rect 1078 148 1097 151
rect 1202 148 1209 151
rect 1366 148 1385 151
rect 1414 148 1430 151
rect 1518 148 1526 151
rect 1586 148 1593 151
rect 634 138 641 141
rect 698 138 705 141
rect 930 138 937 141
rect 94 128 113 131
rect 142 131 146 136
rect 142 128 158 131
rect 418 128 419 132
rect 446 128 449 138
rect 478 131 482 136
rect 478 128 494 131
rect 566 128 585 131
rect 702 128 705 138
rect 710 128 729 131
rect 1350 131 1354 133
rect 1350 128 1361 131
rect 29 118 30 122
rect 1170 118 1171 122
rect 1234 118 1235 122
rect 888 103 890 107
rect 894 103 897 107
rect 901 103 904 107
rect 1069 88 1070 92
rect 1370 88 1371 92
rect 222 71 225 81
rect 454 78 465 81
rect 470 78 489 81
rect 838 78 849 81
rect 454 77 458 78
rect 838 77 842 78
rect 222 68 241 71
rect 742 68 754 71
rect 866 68 873 71
rect 1350 71 1354 74
rect 1350 68 1358 71
rect 1402 68 1425 71
rect 1494 68 1502 71
rect 398 58 414 61
rect 854 58 873 61
rect 930 58 937 61
rect 1118 58 1126 61
rect 1206 58 1214 61
rect 1238 58 1249 61
rect 1390 58 1425 61
rect 1454 58 1462 61
rect 1062 42 1066 44
rect 368 3 370 7
rect 374 3 377 7
rect 381 3 384 7
rect 1384 3 1386 7
rect 1390 3 1393 7
rect 1397 3 1400 7
<< m2contact >>
rect 890 1703 894 1707
rect 897 1703 901 1707
rect 158 1688 162 1692
rect 526 1688 530 1692
rect 1550 1688 1554 1692
rect 1766 1688 1770 1692
rect 14 1678 18 1682
rect 430 1678 434 1682
rect 1254 1678 1258 1682
rect 1438 1678 1442 1682
rect 342 1668 346 1672
rect 414 1668 418 1672
rect 598 1668 602 1672
rect 614 1668 618 1672
rect 702 1668 706 1672
rect 742 1668 746 1672
rect 814 1668 818 1672
rect 854 1668 858 1672
rect 918 1668 922 1672
rect 1046 1668 1050 1672
rect 1126 1668 1130 1672
rect 1270 1668 1274 1672
rect 1422 1668 1426 1672
rect 1566 1668 1570 1672
rect 54 1658 58 1662
rect 62 1658 66 1662
rect 94 1659 98 1663
rect 126 1658 130 1662
rect 206 1658 210 1662
rect 222 1658 226 1662
rect 326 1659 330 1663
rect 374 1658 378 1662
rect 382 1658 386 1662
rect 462 1659 466 1663
rect 494 1658 498 1662
rect 534 1658 538 1662
rect 638 1658 642 1662
rect 806 1658 810 1662
rect 886 1658 890 1662
rect 942 1658 946 1662
rect 1006 1658 1010 1662
rect 1014 1658 1018 1662
rect 1118 1658 1122 1662
rect 1302 1658 1306 1662
rect 1318 1658 1322 1662
rect 1478 1658 1482 1662
rect 1590 1658 1594 1662
rect 1654 1658 1658 1662
rect 1662 1658 1666 1662
rect 1686 1658 1690 1662
rect 1702 1658 1706 1662
rect 1710 1658 1714 1662
rect 1734 1658 1738 1662
rect 1742 1658 1746 1662
rect 1774 1658 1778 1662
rect 38 1648 42 1652
rect 1318 1648 1322 1652
rect 1366 1648 1370 1652
rect 1390 1650 1394 1654
rect 678 1638 682 1642
rect 1390 1627 1394 1631
rect 254 1618 258 1622
rect 262 1618 266 1622
rect 694 1618 698 1622
rect 726 1618 730 1622
rect 838 1618 842 1622
rect 998 1618 1002 1622
rect 1070 1618 1074 1622
rect 1174 1618 1178 1622
rect 1318 1618 1322 1622
rect 1518 1618 1522 1622
rect 1646 1618 1650 1622
rect 1678 1618 1682 1622
rect 1726 1618 1730 1622
rect 1790 1618 1794 1622
rect 370 1603 374 1607
rect 377 1603 381 1607
rect 1386 1603 1390 1607
rect 1393 1603 1397 1607
rect 206 1588 210 1592
rect 286 1588 290 1592
rect 926 1588 930 1592
rect 1750 1588 1754 1592
rect 1798 1588 1802 1592
rect 534 1578 538 1582
rect 1590 1579 1594 1583
rect 102 1568 106 1572
rect 1014 1568 1018 1572
rect 1150 1568 1154 1572
rect 182 1558 186 1562
rect 270 1558 274 1562
rect 598 1558 602 1562
rect 1590 1556 1594 1560
rect 38 1548 42 1552
rect 62 1548 66 1552
rect 150 1548 154 1552
rect 158 1548 162 1552
rect 190 1548 194 1552
rect 198 1548 202 1552
rect 398 1548 402 1552
rect 422 1548 426 1552
rect 478 1548 482 1552
rect 510 1548 514 1552
rect 518 1548 522 1552
rect 526 1548 530 1552
rect 606 1548 610 1552
rect 614 1548 618 1552
rect 702 1548 706 1552
rect 726 1548 730 1552
rect 766 1548 770 1552
rect 822 1547 826 1551
rect 910 1548 914 1552
rect 918 1548 922 1552
rect 1022 1548 1026 1552
rect 1030 1548 1034 1552
rect 1094 1548 1098 1552
rect 1190 1548 1194 1552
rect 1278 1548 1282 1552
rect 1286 1548 1290 1552
rect 1294 1548 1298 1552
rect 1302 1548 1306 1552
rect 1398 1547 1402 1551
rect 1574 1548 1578 1552
rect 1734 1548 1738 1552
rect 1774 1548 1778 1552
rect 118 1538 122 1542
rect 166 1538 170 1542
rect 254 1538 258 1542
rect 342 1538 346 1542
rect 358 1538 362 1542
rect 502 1538 506 1542
rect 574 1538 578 1542
rect 646 1538 650 1542
rect 750 1538 754 1542
rect 774 1538 778 1542
rect 790 1538 794 1542
rect 806 1538 810 1542
rect 1190 1538 1194 1542
rect 1254 1538 1258 1542
rect 1334 1538 1338 1542
rect 1470 1538 1474 1542
rect 1622 1538 1626 1542
rect 102 1528 106 1532
rect 686 1528 690 1532
rect 790 1528 794 1532
rect 966 1528 970 1532
rect 974 1528 978 1532
rect 1102 1528 1106 1532
rect 1230 1528 1234 1532
rect 1350 1528 1354 1532
rect 1398 1528 1402 1532
rect 1542 1528 1546 1532
rect 1638 1528 1642 1532
rect 1766 1528 1770 1532
rect 182 1518 186 1522
rect 270 1518 274 1522
rect 454 1518 458 1522
rect 494 1518 498 1522
rect 590 1518 594 1522
rect 886 1518 890 1522
rect 1038 1518 1042 1522
rect 1134 1518 1138 1522
rect 1462 1518 1466 1522
rect 1526 1518 1530 1522
rect 1550 1518 1554 1522
rect 1718 1518 1722 1522
rect 1758 1518 1762 1522
rect 890 1503 894 1507
rect 897 1503 901 1507
rect 94 1488 98 1492
rect 558 1488 562 1492
rect 678 1488 682 1492
rect 790 1488 794 1492
rect 1014 1488 1018 1492
rect 1118 1488 1122 1492
rect 1502 1488 1506 1492
rect 1582 1488 1586 1492
rect 102 1478 106 1482
rect 206 1478 210 1482
rect 438 1478 442 1482
rect 494 1478 498 1482
rect 630 1478 634 1482
rect 750 1478 754 1482
rect 798 1478 802 1482
rect 990 1478 994 1482
rect 1086 1478 1090 1482
rect 126 1468 130 1472
rect 142 1468 146 1472
rect 158 1468 162 1472
rect 254 1468 258 1472
rect 358 1468 362 1472
rect 398 1468 402 1472
rect 446 1468 450 1472
rect 598 1468 602 1472
rect 638 1468 642 1472
rect 670 1468 674 1472
rect 846 1468 850 1472
rect 934 1468 938 1472
rect 998 1468 1002 1472
rect 1014 1468 1018 1472
rect 1046 1468 1050 1472
rect 1054 1468 1058 1472
rect 1070 1468 1074 1472
rect 1310 1468 1314 1472
rect 1470 1468 1474 1472
rect 1494 1468 1498 1472
rect 1518 1478 1522 1482
rect 1558 1478 1562 1482
rect 1614 1478 1618 1482
rect 1702 1478 1706 1482
rect 1574 1468 1578 1472
rect 1686 1468 1690 1472
rect 38 1458 42 1462
rect 62 1458 66 1462
rect 118 1458 122 1462
rect 150 1458 154 1462
rect 190 1458 194 1462
rect 214 1458 218 1462
rect 222 1458 226 1462
rect 334 1458 338 1462
rect 390 1458 394 1462
rect 422 1458 426 1462
rect 494 1459 498 1463
rect 574 1458 578 1462
rect 646 1458 650 1462
rect 750 1459 754 1463
rect 782 1458 786 1462
rect 806 1458 810 1462
rect 814 1458 818 1462
rect 942 1458 946 1462
rect 1006 1458 1010 1462
rect 1046 1458 1050 1462
rect 1086 1458 1090 1462
rect 1134 1458 1138 1462
rect 1142 1458 1146 1462
rect 1150 1458 1154 1462
rect 1158 1458 1162 1462
rect 1246 1458 1250 1462
rect 1270 1458 1274 1462
rect 1318 1458 1322 1462
rect 1342 1458 1346 1462
rect 1350 1458 1354 1462
rect 1366 1458 1370 1462
rect 1446 1458 1450 1462
rect 1486 1458 1490 1462
rect 1542 1458 1546 1462
rect 1566 1458 1570 1462
rect 1598 1458 1602 1462
rect 1646 1458 1650 1462
rect 174 1448 178 1452
rect 414 1448 418 1452
rect 462 1448 466 1452
rect 614 1448 618 1452
rect 982 1448 986 1452
rect 1174 1448 1178 1452
rect 1326 1448 1330 1452
rect 1654 1450 1658 1454
rect 182 1438 186 1442
rect 590 1438 594 1442
rect 278 1418 282 1422
rect 454 1418 458 1422
rect 582 1418 586 1422
rect 886 1418 890 1422
rect 1070 1418 1074 1422
rect 1214 1418 1218 1422
rect 1542 1418 1546 1422
rect 1654 1418 1658 1422
rect 1782 1418 1786 1422
rect 370 1403 374 1407
rect 377 1403 381 1407
rect 1386 1403 1390 1407
rect 1393 1403 1397 1407
rect 286 1388 290 1392
rect 574 1388 578 1392
rect 750 1388 754 1392
rect 1630 1388 1634 1392
rect 1742 1388 1746 1392
rect 190 1368 194 1372
rect 262 1368 266 1372
rect 334 1368 338 1372
rect 366 1368 370 1372
rect 566 1368 570 1372
rect 622 1368 626 1372
rect 254 1358 258 1362
rect 310 1358 314 1362
rect 318 1358 322 1362
rect 550 1358 554 1362
rect 598 1358 602 1362
rect 606 1358 610 1362
rect 654 1358 658 1362
rect 662 1358 666 1362
rect 702 1358 706 1362
rect 774 1358 778 1362
rect 798 1358 802 1362
rect 918 1358 922 1362
rect 1486 1358 1490 1362
rect 1638 1358 1642 1362
rect 1782 1358 1786 1362
rect 30 1347 34 1351
rect 62 1348 66 1352
rect 134 1348 138 1352
rect 198 1348 202 1352
rect 206 1348 210 1352
rect 222 1348 226 1352
rect 270 1348 274 1352
rect 310 1348 314 1352
rect 326 1348 330 1352
rect 358 1348 362 1352
rect 438 1348 442 1352
rect 494 1348 498 1352
rect 542 1348 546 1352
rect 558 1348 562 1352
rect 614 1348 618 1352
rect 718 1348 722 1352
rect 726 1348 730 1352
rect 734 1348 738 1352
rect 758 1348 762 1352
rect 846 1348 850 1352
rect 878 1348 882 1352
rect 926 1348 930 1352
rect 958 1348 962 1352
rect 110 1338 114 1342
rect 158 1338 162 1342
rect 294 1338 298 1342
rect 1030 1347 1034 1351
rect 1062 1348 1066 1352
rect 1078 1348 1082 1352
rect 1102 1348 1106 1352
rect 1150 1348 1154 1352
rect 1158 1348 1162 1352
rect 1198 1348 1202 1352
rect 1262 1348 1266 1352
rect 1278 1348 1282 1352
rect 1310 1348 1314 1352
rect 1318 1348 1322 1352
rect 1326 1348 1330 1352
rect 1342 1348 1346 1352
rect 1358 1348 1362 1352
rect 1374 1348 1378 1352
rect 1446 1348 1450 1352
rect 1566 1348 1570 1352
rect 1574 1348 1578 1352
rect 1606 1348 1610 1352
rect 1630 1348 1634 1352
rect 1662 1348 1666 1352
rect 1678 1348 1682 1352
rect 1686 1348 1690 1352
rect 1710 1348 1714 1352
rect 1726 1348 1730 1352
rect 1734 1348 1738 1352
rect 1758 1348 1762 1352
rect 430 1338 434 1342
rect 526 1338 530 1342
rect 534 1338 538 1342
rect 582 1338 586 1342
rect 638 1338 642 1342
rect 678 1338 682 1342
rect 686 1338 690 1342
rect 790 1338 794 1342
rect 814 1338 818 1342
rect 838 1338 842 1342
rect 878 1338 882 1342
rect 934 1338 938 1342
rect 950 1338 954 1342
rect 1030 1338 1034 1342
rect 1070 1338 1074 1342
rect 1086 1338 1090 1342
rect 1190 1338 1194 1342
rect 1278 1338 1282 1342
rect 1470 1338 1474 1342
rect 1510 1338 1514 1342
rect 1598 1338 1602 1342
rect 1670 1338 1674 1342
rect 1782 1338 1786 1342
rect 254 1328 258 1332
rect 382 1328 386 1332
rect 510 1328 514 1332
rect 718 1328 722 1332
rect 830 1328 834 1332
rect 1102 1328 1106 1332
rect 1518 1328 1522 1332
rect 1598 1328 1602 1332
rect 1798 1328 1802 1332
rect 94 1318 98 1322
rect 486 1318 490 1322
rect 598 1318 602 1322
rect 622 1318 626 1322
rect 646 1318 650 1322
rect 670 1318 674 1322
rect 702 1318 706 1322
rect 774 1318 778 1322
rect 806 1318 810 1322
rect 886 1318 890 1322
rect 942 1318 946 1322
rect 966 1318 970 1322
rect 1134 1318 1138 1322
rect 1390 1318 1394 1322
rect 1486 1318 1490 1322
rect 1550 1318 1554 1322
rect 1694 1318 1698 1322
rect 890 1303 894 1307
rect 897 1303 901 1307
rect 30 1288 34 1292
rect 222 1288 226 1292
rect 350 1288 354 1292
rect 590 1288 594 1292
rect 798 1288 802 1292
rect 1038 1288 1042 1292
rect 1078 1288 1082 1292
rect 1174 1288 1178 1292
rect 1422 1288 1426 1292
rect 1478 1288 1482 1292
rect 1502 1288 1506 1292
rect 62 1278 66 1282
rect 126 1278 130 1282
rect 158 1278 162 1282
rect 390 1278 394 1282
rect 430 1278 434 1282
rect 454 1278 458 1282
rect 494 1278 498 1282
rect 526 1278 530 1282
rect 606 1278 610 1282
rect 758 1278 762 1282
rect 1070 1278 1074 1282
rect 1206 1278 1210 1282
rect 1238 1278 1242 1282
rect 1270 1278 1274 1282
rect 1302 1278 1306 1282
rect 1390 1278 1394 1282
rect 1430 1278 1434 1282
rect 1494 1278 1498 1282
rect 1702 1278 1706 1282
rect 110 1268 114 1272
rect 126 1268 130 1272
rect 270 1268 274 1272
rect 510 1268 514 1272
rect 766 1268 770 1272
rect 854 1268 858 1272
rect 950 1268 954 1272
rect 998 1268 1002 1272
rect 1014 1268 1018 1272
rect 1030 1268 1034 1272
rect 1158 1268 1162 1272
rect 1270 1268 1274 1272
rect 1334 1268 1338 1272
rect 1350 1268 1354 1272
rect 1366 1268 1370 1272
rect 1406 1268 1410 1272
rect 1486 1268 1490 1272
rect 1558 1268 1562 1272
rect 1598 1268 1602 1272
rect 1614 1268 1618 1272
rect 1630 1268 1634 1272
rect 1750 1268 1754 1272
rect 14 1258 18 1262
rect 38 1258 42 1262
rect 46 1258 50 1262
rect 62 1258 66 1262
rect 70 1258 74 1262
rect 78 1258 82 1262
rect 158 1259 162 1263
rect 238 1258 242 1262
rect 294 1258 298 1262
rect 374 1258 378 1262
rect 382 1258 386 1262
rect 438 1258 442 1262
rect 446 1258 450 1262
rect 534 1258 538 1262
rect 614 1258 618 1262
rect 638 1258 642 1262
rect 654 1258 658 1262
rect 678 1258 682 1262
rect 702 1258 706 1262
rect 734 1258 738 1262
rect 782 1258 786 1262
rect 862 1258 866 1262
rect 982 1258 986 1262
rect 990 1258 994 1262
rect 1022 1258 1026 1262
rect 1054 1258 1058 1262
rect 1134 1258 1138 1262
rect 1238 1259 1242 1263
rect 1286 1258 1290 1262
rect 1294 1258 1298 1262
rect 1318 1258 1322 1262
rect 1342 1258 1346 1262
rect 1358 1258 1362 1262
rect 1406 1258 1410 1262
rect 1470 1258 1474 1262
rect 1534 1258 1538 1262
rect 1550 1258 1554 1262
rect 1606 1258 1610 1262
rect 1622 1258 1626 1262
rect 1630 1258 1634 1262
rect 1646 1258 1650 1262
rect 1670 1258 1674 1262
rect 1686 1258 1690 1262
rect 1734 1259 1738 1263
rect 1766 1258 1770 1262
rect 206 1248 210 1252
rect 230 1248 234 1252
rect 622 1248 626 1252
rect 630 1248 634 1252
rect 686 1248 690 1252
rect 246 1238 250 1242
rect 606 1238 610 1242
rect 646 1238 650 1242
rect 670 1238 674 1242
rect 726 1248 730 1252
rect 998 1248 1002 1252
rect 1662 1248 1666 1252
rect 710 1238 714 1242
rect 742 1238 746 1242
rect 934 1238 938 1242
rect 254 1218 258 1222
rect 718 1218 722 1222
rect 750 1218 754 1222
rect 1686 1218 1690 1222
rect 1798 1218 1802 1222
rect 370 1203 374 1207
rect 377 1203 381 1207
rect 1386 1203 1390 1207
rect 1393 1203 1397 1207
rect 398 1188 402 1192
rect 814 1188 818 1192
rect 958 1178 962 1182
rect 1606 1178 1610 1182
rect 30 1168 34 1172
rect 158 1168 162 1172
rect 438 1168 442 1172
rect 566 1168 570 1172
rect 806 1168 810 1172
rect 998 1168 1002 1172
rect 1390 1168 1394 1172
rect 406 1158 410 1162
rect 550 1158 554 1162
rect 814 1158 818 1162
rect 830 1158 834 1162
rect 974 1158 978 1162
rect 1126 1158 1130 1162
rect 1694 1158 1698 1162
rect 1726 1158 1730 1162
rect 14 1148 18 1152
rect 38 1148 42 1152
rect 46 1148 50 1152
rect 62 1148 66 1152
rect 94 1147 98 1151
rect 126 1148 130 1152
rect 166 1148 170 1152
rect 198 1148 202 1152
rect 254 1148 258 1152
rect 270 1148 274 1152
rect 318 1148 322 1152
rect 350 1148 354 1152
rect 414 1148 418 1152
rect 422 1148 426 1152
rect 502 1147 506 1151
rect 630 1148 634 1152
rect 718 1148 722 1152
rect 726 1148 730 1152
rect 758 1148 762 1152
rect 814 1148 818 1152
rect 854 1148 858 1152
rect 862 1148 866 1152
rect 926 1148 930 1152
rect 966 1148 970 1152
rect 1054 1148 1058 1152
rect 1142 1148 1146 1152
rect 1150 1148 1154 1152
rect 1214 1148 1218 1152
rect 1326 1148 1330 1152
rect 1334 1148 1338 1152
rect 1438 1148 1442 1152
rect 1462 1148 1466 1152
rect 1550 1148 1554 1152
rect 1614 1148 1618 1152
rect 1622 1148 1626 1152
rect 1710 1148 1714 1152
rect 1734 1148 1738 1152
rect 174 1138 178 1142
rect 326 1138 330 1142
rect 366 1138 370 1142
rect 510 1138 514 1142
rect 654 1138 658 1142
rect 734 1138 738 1142
rect 830 1138 834 1142
rect 846 1138 850 1142
rect 910 1138 914 1142
rect 934 1138 938 1142
rect 958 1138 962 1142
rect 990 1138 994 1142
rect 1054 1138 1058 1142
rect 1078 1138 1082 1142
rect 1214 1138 1218 1142
rect 1318 1138 1322 1142
rect 1366 1138 1370 1142
rect 1526 1138 1530 1142
rect 1670 1138 1674 1142
rect 1702 1138 1706 1142
rect 62 1128 66 1132
rect 214 1128 218 1132
rect 246 1128 250 1132
rect 334 1128 338 1132
rect 366 1128 370 1132
rect 470 1128 474 1132
rect 670 1128 674 1132
rect 742 1128 746 1132
rect 926 1128 930 1132
rect 1094 1128 1098 1132
rect 1510 1128 1514 1132
rect 1630 1128 1634 1132
rect 1742 1128 1746 1132
rect 182 1118 186 1122
rect 310 1118 314 1122
rect 574 1118 578 1122
rect 710 1118 714 1122
rect 790 1118 794 1122
rect 974 1118 978 1122
rect 1158 1118 1162 1122
rect 1262 1118 1266 1122
rect 1502 1118 1506 1122
rect 1686 1118 1690 1122
rect 1750 1118 1754 1122
rect 890 1103 894 1107
rect 897 1103 901 1107
rect 382 1088 386 1092
rect 510 1088 514 1092
rect 542 1088 546 1092
rect 598 1088 602 1092
rect 678 1088 682 1092
rect 854 1088 858 1092
rect 878 1088 882 1092
rect 1038 1088 1042 1092
rect 1070 1088 1074 1092
rect 1110 1088 1114 1092
rect 1614 1088 1618 1092
rect 1646 1088 1650 1092
rect 1678 1088 1682 1092
rect 150 1078 154 1082
rect 214 1078 218 1082
rect 462 1078 466 1082
rect 582 1078 586 1082
rect 110 1068 114 1072
rect 166 1068 170 1072
rect 262 1068 266 1072
rect 278 1068 282 1072
rect 302 1068 306 1072
rect 470 1068 474 1072
rect 534 1068 538 1072
rect 550 1068 554 1072
rect 782 1078 786 1082
rect 822 1078 826 1082
rect 1094 1078 1098 1082
rect 1478 1078 1482 1082
rect 1558 1078 1562 1082
rect 1686 1078 1690 1082
rect 606 1068 610 1072
rect 654 1068 658 1072
rect 670 1068 674 1072
rect 758 1068 762 1072
rect 782 1068 786 1072
rect 830 1068 834 1072
rect 862 1068 866 1072
rect 910 1068 914 1072
rect 982 1068 986 1072
rect 998 1068 1002 1072
rect 1014 1068 1018 1072
rect 1030 1068 1034 1072
rect 1062 1068 1066 1072
rect 1078 1068 1082 1072
rect 1214 1068 1218 1072
rect 1310 1068 1314 1072
rect 1358 1068 1362 1072
rect 1438 1068 1442 1072
rect 1590 1068 1594 1072
rect 1622 1068 1626 1072
rect 1654 1068 1658 1072
rect 1670 1068 1674 1072
rect 1766 1068 1770 1072
rect 38 1058 42 1062
rect 62 1058 66 1062
rect 102 1058 106 1062
rect 118 1058 122 1062
rect 134 1058 138 1062
rect 182 1059 186 1063
rect 286 1058 290 1062
rect 326 1058 330 1062
rect 398 1058 402 1062
rect 414 1058 418 1062
rect 502 1058 506 1062
rect 526 1058 530 1062
rect 558 1058 562 1062
rect 566 1058 570 1062
rect 614 1058 618 1062
rect 630 1058 634 1062
rect 718 1058 722 1062
rect 798 1058 802 1062
rect 822 1058 826 1062
rect 870 1058 874 1062
rect 990 1058 994 1062
rect 1006 1058 1010 1062
rect 1022 1058 1026 1062
rect 1046 1058 1050 1062
rect 1094 1058 1098 1062
rect 1166 1058 1170 1062
rect 1230 1059 1234 1063
rect 1262 1058 1266 1062
rect 1342 1058 1346 1062
rect 1430 1058 1434 1062
rect 1438 1058 1442 1062
rect 1462 1058 1466 1062
rect 1470 1058 1474 1062
rect 1478 1058 1482 1062
rect 1558 1059 1562 1063
rect 1598 1058 1602 1062
rect 1630 1058 1634 1062
rect 1646 1058 1650 1062
rect 1662 1058 1666 1062
rect 1702 1058 1706 1062
rect 1766 1058 1770 1062
rect 430 1048 434 1052
rect 470 1048 474 1052
rect 486 1048 490 1052
rect 518 1048 522 1052
rect 622 1048 626 1052
rect 654 1048 658 1052
rect 878 1048 882 1052
rect 1614 1048 1618 1052
rect 502 1038 506 1042
rect 638 1038 642 1042
rect 694 1038 698 1042
rect 1494 1038 1498 1042
rect 1726 1038 1730 1042
rect 278 1028 282 1032
rect 94 1018 98 1022
rect 630 1018 634 1022
rect 926 1018 930 1022
rect 1038 1018 1042 1022
rect 1102 1018 1106 1022
rect 1294 1018 1298 1022
rect 370 1003 374 1007
rect 377 1003 381 1007
rect 1386 1003 1390 1007
rect 1393 1003 1397 1007
rect 454 988 458 992
rect 478 988 482 992
rect 510 988 514 992
rect 678 988 682 992
rect 862 988 866 992
rect 966 988 970 992
rect 1006 988 1010 992
rect 1126 988 1130 992
rect 1382 988 1386 992
rect 1558 988 1562 992
rect 1766 988 1770 992
rect 1790 988 1794 992
rect 1310 979 1314 983
rect 94 968 98 972
rect 374 968 378 972
rect 446 968 450 972
rect 486 968 490 972
rect 766 968 770 972
rect 358 958 362 962
rect 462 958 466 962
rect 470 958 474 962
rect 502 958 506 962
rect 974 958 978 962
rect 998 958 1002 962
rect 1310 956 1314 960
rect 1382 958 1386 962
rect 1606 958 1610 962
rect 38 948 42 952
rect 150 948 154 952
rect 158 948 162 952
rect 166 948 170 952
rect 198 948 202 952
rect 206 948 210 952
rect 238 948 242 952
rect 254 948 258 952
rect 302 948 306 952
rect 366 948 370 952
rect 414 948 418 952
rect 454 948 458 952
rect 478 948 482 952
rect 574 948 578 952
rect 622 948 626 952
rect 646 948 650 952
rect 734 948 738 952
rect 742 948 746 952
rect 806 948 810 952
rect 910 948 914 952
rect 1046 948 1050 952
rect 1102 948 1106 952
rect 1134 948 1138 952
rect 1142 948 1146 952
rect 1150 948 1154 952
rect 1326 948 1330 952
rect 1374 948 1378 952
rect 1486 948 1490 952
rect 1550 948 1554 952
rect 1574 948 1578 952
rect 1582 948 1586 952
rect 1598 948 1602 952
rect 1622 948 1626 952
rect 1630 948 1634 952
rect 1646 948 1650 952
rect 1710 948 1714 952
rect 1750 948 1754 952
rect 1774 948 1778 952
rect 118 938 122 942
rect 174 938 178 942
rect 206 938 210 942
rect 246 938 250 942
rect 310 938 314 942
rect 406 938 410 942
rect 518 938 522 942
rect 566 938 570 942
rect 598 938 602 942
rect 702 938 706 942
rect 830 938 834 942
rect 926 938 930 942
rect 958 938 962 942
rect 982 938 986 942
rect 1054 938 1058 942
rect 1062 938 1066 942
rect 1278 938 1282 942
rect 1430 938 1434 942
rect 1734 938 1738 942
rect 30 928 34 932
rect 222 928 226 932
rect 574 928 578 932
rect 1150 928 1154 932
rect 1182 928 1186 932
rect 1262 928 1266 932
rect 1446 928 1450 932
rect 190 918 194 922
rect 262 918 266 922
rect 366 918 370 922
rect 430 918 434 922
rect 566 918 570 922
rect 750 918 754 922
rect 854 918 858 922
rect 998 918 1002 922
rect 1526 918 1530 922
rect 890 903 894 907
rect 897 903 901 907
rect 94 888 98 892
rect 182 888 186 892
rect 422 888 426 892
rect 454 888 458 892
rect 470 888 474 892
rect 582 888 586 892
rect 646 888 650 892
rect 734 888 738 892
rect 846 888 850 892
rect 910 888 914 892
rect 966 888 970 892
rect 1158 888 1162 892
rect 1206 888 1210 892
rect 1358 888 1362 892
rect 1606 888 1610 892
rect 1734 888 1738 892
rect 1798 888 1802 892
rect 30 878 34 882
rect 102 878 106 882
rect 134 878 138 882
rect 150 878 154 882
rect 254 878 258 882
rect 302 878 306 882
rect 102 868 106 872
rect 118 868 122 872
rect 174 868 178 872
rect 206 868 210 872
rect 214 868 218 872
rect 294 868 298 872
rect 38 858 42 862
rect 62 858 66 862
rect 126 858 130 862
rect 198 858 202 862
rect 254 858 258 862
rect 286 858 290 862
rect 390 868 394 872
rect 430 868 434 872
rect 446 868 450 872
rect 550 868 554 872
rect 574 868 578 872
rect 598 878 602 882
rect 702 878 706 882
rect 854 878 858 882
rect 934 878 938 882
rect 1014 878 1018 882
rect 1062 878 1066 882
rect 1150 878 1154 882
rect 1238 878 1242 882
rect 1270 878 1274 882
rect 1406 878 1410 882
rect 1494 878 1498 882
rect 1574 878 1578 882
rect 1670 878 1674 882
rect 1734 878 1738 882
rect 622 868 626 872
rect 678 868 682 872
rect 694 868 698 872
rect 742 868 746 872
rect 798 868 802 872
rect 822 868 826 872
rect 830 868 834 872
rect 990 868 994 872
rect 1166 868 1170 872
rect 1350 868 1354 872
rect 1478 868 1482 872
rect 1598 868 1602 872
rect 1638 868 1642 872
rect 1646 868 1650 872
rect 1678 868 1682 872
rect 1686 868 1690 872
rect 318 858 322 862
rect 342 855 346 859
rect 374 858 378 862
rect 406 858 410 862
rect 438 858 442 862
rect 534 859 538 863
rect 566 858 570 862
rect 614 858 618 862
rect 662 858 666 862
rect 718 858 722 862
rect 750 858 754 862
rect 758 858 762 862
rect 766 858 770 862
rect 790 858 794 862
rect 918 858 922 862
rect 934 858 938 862
rect 950 858 954 862
rect 982 858 986 862
rect 998 858 1002 862
rect 1022 858 1026 862
rect 1030 858 1034 862
rect 1062 859 1066 863
rect 1174 858 1178 862
rect 1190 858 1194 862
rect 1214 858 1218 862
rect 1222 858 1226 862
rect 1278 858 1282 862
rect 1342 858 1346 862
rect 1374 858 1378 862
rect 1534 858 1538 862
rect 1590 858 1594 862
rect 1622 858 1626 862
rect 1654 858 1658 862
rect 1670 858 1674 862
rect 1694 858 1698 862
rect 1710 858 1714 862
rect 1782 858 1786 862
rect 174 848 178 852
rect 230 848 234 852
rect 262 848 266 852
rect 270 848 274 852
rect 350 848 354 852
rect 462 848 466 852
rect 638 848 642 852
rect 678 848 682 852
rect 694 848 698 852
rect 806 848 810 852
rect 846 848 850 852
rect 1238 848 1242 852
rect 1446 850 1450 854
rect 1710 848 1714 852
rect 246 838 250 842
rect 366 838 370 842
rect 654 838 658 842
rect 182 818 186 822
rect 222 818 226 822
rect 278 818 282 822
rect 390 818 394 822
rect 630 818 634 822
rect 782 818 786 822
rect 1142 818 1146 822
rect 1334 818 1338 822
rect 1446 818 1450 822
rect 370 803 374 807
rect 377 803 381 807
rect 1386 803 1390 807
rect 1393 803 1397 807
rect 214 788 218 792
rect 254 788 258 792
rect 350 788 354 792
rect 446 788 450 792
rect 742 788 746 792
rect 790 788 794 792
rect 966 788 970 792
rect 1006 788 1010 792
rect 1158 788 1162 792
rect 1334 788 1338 792
rect 1702 788 1706 792
rect 1134 778 1138 782
rect 1510 779 1514 783
rect 126 768 130 772
rect 230 768 234 772
rect 246 768 250 772
rect 574 768 578 772
rect 766 768 770 772
rect 1230 768 1234 772
rect 1382 768 1386 772
rect 134 758 138 762
rect 222 758 226 762
rect 230 758 234 762
rect 454 758 458 762
rect 558 758 562 762
rect 974 758 978 762
rect 1126 758 1130 762
rect 1510 756 1514 760
rect 38 748 42 752
rect 62 748 66 752
rect 190 748 194 752
rect 198 748 202 752
rect 238 748 242 752
rect 294 748 298 752
rect 318 748 322 752
rect 422 748 426 752
rect 430 748 434 752
rect 494 748 498 752
rect 614 748 618 752
rect 630 748 634 752
rect 726 748 730 752
rect 734 748 738 752
rect 758 748 762 752
rect 766 748 770 752
rect 806 748 810 752
rect 822 748 826 752
rect 838 748 842 752
rect 910 748 914 752
rect 1006 748 1010 752
rect 1046 748 1050 752
rect 1054 748 1058 752
rect 1062 748 1066 752
rect 1086 748 1090 752
rect 1110 748 1114 752
rect 1182 748 1186 752
rect 1222 748 1226 752
rect 1238 748 1242 752
rect 1254 748 1258 752
rect 1262 748 1266 752
rect 1286 748 1290 752
rect 1326 748 1330 752
rect 1350 748 1354 752
rect 1358 748 1362 752
rect 1374 748 1378 752
rect 1438 748 1442 752
rect 1542 748 1546 752
rect 1654 748 1658 752
rect 1662 748 1666 752
rect 1694 748 1698 752
rect 1758 748 1762 752
rect 158 738 162 742
rect 206 738 210 742
rect 374 738 378 742
rect 438 738 442 742
rect 470 738 474 742
rect 574 738 578 742
rect 702 738 706 742
rect 782 738 786 742
rect 814 738 818 742
rect 830 738 834 742
rect 926 738 930 742
rect 958 738 962 742
rect 982 738 986 742
rect 1006 738 1010 742
rect 1102 738 1106 742
rect 1126 738 1130 742
rect 1142 738 1146 742
rect 1158 738 1162 742
rect 1182 738 1186 742
rect 1214 738 1218 742
rect 1246 738 1250 742
rect 1294 738 1298 742
rect 1542 738 1546 742
rect 1686 738 1690 742
rect 1758 738 1762 742
rect 110 728 114 732
rect 142 728 146 732
rect 646 728 650 732
rect 678 728 682 732
rect 1030 728 1034 732
rect 1046 728 1050 732
rect 1158 728 1162 732
rect 1190 728 1194 732
rect 1310 728 1314 732
rect 1446 728 1450 732
rect 1558 728 1562 732
rect 94 718 98 722
rect 102 718 106 722
rect 550 718 554 722
rect 558 718 562 722
rect 862 718 866 722
rect 974 718 978 722
rect 1014 718 1018 722
rect 1078 718 1082 722
rect 1638 718 1642 722
rect 890 703 894 707
rect 897 703 901 707
rect 94 688 98 692
rect 238 688 242 692
rect 278 688 282 692
rect 390 688 394 692
rect 638 688 642 692
rect 670 688 674 692
rect 694 688 698 692
rect 790 688 794 692
rect 870 688 874 692
rect 910 688 914 692
rect 1166 688 1170 692
rect 1182 688 1186 692
rect 1470 688 1474 692
rect 1534 688 1538 692
rect 1798 688 1802 692
rect 270 678 274 682
rect 6 668 10 672
rect 78 668 82 672
rect 158 668 162 672
rect 238 668 242 672
rect 254 668 258 672
rect 270 668 274 672
rect 382 668 386 672
rect 470 668 474 672
rect 486 668 490 672
rect 502 668 506 672
rect 518 678 522 682
rect 550 678 554 682
rect 598 678 602 682
rect 726 678 730 682
rect 982 678 986 682
rect 1014 678 1018 682
rect 1102 678 1106 682
rect 1174 678 1178 682
rect 1270 678 1274 682
rect 1462 678 1466 682
rect 1542 678 1546 682
rect 1670 678 1674 682
rect 1686 678 1690 682
rect 1758 678 1762 682
rect 1790 678 1794 682
rect 542 668 546 672
rect 646 668 650 672
rect 678 668 682 672
rect 686 668 690 672
rect 814 668 818 672
rect 862 668 866 672
rect 910 668 914 672
rect 1030 668 1034 672
rect 1230 668 1234 672
rect 1358 668 1362 672
rect 1390 668 1394 672
rect 1414 668 1418 672
rect 1446 668 1450 672
rect 1478 668 1482 672
rect 1502 668 1506 672
rect 1518 668 1522 672
rect 1526 668 1530 672
rect 1542 668 1546 672
rect 1574 668 1578 672
rect 1630 668 1634 672
rect 1662 668 1666 672
rect 1742 668 1746 672
rect 46 658 50 662
rect 54 658 58 662
rect 86 658 90 662
rect 150 658 154 662
rect 190 658 194 662
rect 198 658 202 662
rect 222 658 226 662
rect 318 658 322 662
rect 334 658 338 662
rect 422 658 426 662
rect 454 659 458 663
rect 486 658 490 662
rect 534 658 538 662
rect 566 658 570 662
rect 598 658 602 662
rect 622 658 626 662
rect 662 658 666 662
rect 734 658 738 662
rect 846 658 850 662
rect 854 658 858 662
rect 862 658 866 662
rect 894 658 898 662
rect 982 659 986 663
rect 1062 658 1066 662
rect 1070 658 1074 662
rect 1110 658 1114 662
rect 1190 658 1194 662
rect 1198 658 1202 662
rect 1206 658 1210 662
rect 1238 658 1242 662
rect 1270 659 1274 663
rect 1342 658 1346 662
rect 1366 658 1370 662
rect 1382 658 1386 662
rect 1422 658 1426 662
rect 1438 658 1442 662
rect 1478 658 1482 662
rect 1518 658 1522 662
rect 1582 658 1586 662
rect 1614 658 1618 662
rect 1622 658 1626 662
rect 1638 658 1642 662
rect 1654 658 1658 662
rect 1670 658 1674 662
rect 1734 658 1738 662
rect 238 648 242 652
rect 1438 648 1442 652
rect 1550 648 1554 652
rect 30 618 34 622
rect 1366 618 1370 622
rect 1598 618 1602 622
rect 1638 618 1642 622
rect 1694 618 1698 622
rect 1798 618 1802 622
rect 370 603 374 607
rect 377 603 381 607
rect 1386 603 1390 607
rect 1393 603 1397 607
rect 214 588 218 592
rect 478 588 482 592
rect 526 588 530 592
rect 662 588 666 592
rect 718 588 722 592
rect 822 588 826 592
rect 838 588 842 592
rect 1006 588 1010 592
rect 1174 588 1178 592
rect 1190 588 1194 592
rect 1214 588 1218 592
rect 1678 588 1682 592
rect 1702 588 1706 592
rect 230 568 234 572
rect 406 568 410 572
rect 446 568 450 572
rect 470 568 474 572
rect 566 568 570 572
rect 206 558 210 562
rect 246 558 250 562
rect 278 558 282 562
rect 486 558 490 562
rect 494 558 498 562
rect 1382 558 1386 562
rect 1630 557 1634 561
rect 14 548 18 552
rect 38 548 42 552
rect 46 548 50 552
rect 62 548 66 552
rect 70 548 74 552
rect 102 548 106 552
rect 134 547 138 551
rect 166 548 170 552
rect 254 548 258 552
rect 286 548 290 552
rect 334 547 338 551
rect 406 548 410 552
rect 454 548 458 552
rect 478 548 482 552
rect 558 548 562 552
rect 622 548 626 552
rect 662 548 666 552
rect 702 548 706 552
rect 734 548 738 552
rect 742 548 746 552
rect 790 548 794 552
rect 830 548 834 552
rect 902 547 906 551
rect 950 548 954 552
rect 998 548 1002 552
rect 1070 547 1074 551
rect 1150 548 1154 552
rect 1158 548 1162 552
rect 1238 548 1242 552
rect 1334 547 1338 551
rect 1406 548 1410 552
rect 1430 548 1434 552
rect 1438 548 1442 552
rect 1478 548 1482 552
rect 1542 548 1546 552
rect 1550 548 1554 552
rect 1574 548 1578 552
rect 1614 548 1618 552
rect 1654 548 1658 552
rect 1662 548 1666 552
rect 1686 548 1690 552
rect 1742 548 1746 552
rect 1766 547 1770 551
rect 78 538 82 542
rect 94 538 98 542
rect 222 538 226 542
rect 262 538 266 542
rect 318 538 322 542
rect 366 538 370 542
rect 430 538 434 542
rect 446 538 450 542
rect 494 538 498 542
rect 518 538 522 542
rect 534 538 538 542
rect 614 538 618 542
rect 686 538 690 542
rect 798 538 802 542
rect 822 538 826 542
rect 886 538 890 542
rect 958 538 962 542
rect 1054 538 1058 542
rect 1118 538 1122 542
rect 1182 538 1186 542
rect 1246 538 1250 542
rect 1350 538 1354 542
rect 1382 538 1386 542
rect 1454 538 1458 542
rect 1502 538 1506 542
rect 1606 538 1610 542
rect 302 528 306 532
rect 542 528 546 532
rect 678 528 682 532
rect 686 528 690 532
rect 726 528 730 532
rect 966 528 970 532
rect 982 528 986 532
rect 1102 528 1106 532
rect 1166 528 1170 532
rect 1262 528 1266 532
rect 1366 528 1370 532
rect 1598 528 1602 532
rect 30 518 34 522
rect 86 518 90 522
rect 198 518 202 522
rect 206 518 210 522
rect 550 518 554 522
rect 750 518 754 522
rect 1270 518 1274 522
rect 1534 518 1538 522
rect 1566 518 1570 522
rect 890 503 894 507
rect 897 503 901 507
rect 94 488 98 492
rect 134 488 138 492
rect 190 488 194 492
rect 214 488 218 492
rect 446 488 450 492
rect 510 488 514 492
rect 534 488 538 492
rect 558 488 562 492
rect 646 488 650 492
rect 686 488 690 492
rect 798 488 802 492
rect 902 488 906 492
rect 1006 488 1010 492
rect 1038 488 1042 492
rect 1086 488 1090 492
rect 1182 488 1186 492
rect 1190 488 1194 492
rect 1262 488 1266 492
rect 1326 488 1330 492
rect 1422 488 1426 492
rect 1558 488 1562 492
rect 1566 488 1570 492
rect 1686 488 1690 492
rect 1694 488 1698 492
rect 102 478 106 482
rect 174 478 178 482
rect 350 478 354 482
rect 526 478 530 482
rect 550 478 554 482
rect 598 478 602 482
rect 702 478 706 482
rect 766 478 770 482
rect 934 478 938 482
rect 974 478 978 482
rect 1078 478 1082 482
rect 1222 478 1226 482
rect 1318 478 1322 482
rect 1406 478 1410 482
rect 1702 478 1706 482
rect 166 468 170 472
rect 174 468 178 472
rect 270 468 274 472
rect 318 468 322 472
rect 366 468 370 472
rect 454 468 458 472
rect 566 468 570 472
rect 582 468 586 472
rect 606 468 610 472
rect 646 468 650 472
rect 670 468 674 472
rect 718 468 722 472
rect 814 468 818 472
rect 990 468 994 472
rect 1006 468 1010 472
rect 1014 468 1018 472
rect 1046 468 1050 472
rect 1062 468 1066 472
rect 1102 468 1106 472
rect 1214 468 1218 472
rect 1238 468 1242 472
rect 1270 468 1274 472
rect 1478 468 1482 472
rect 1534 468 1538 472
rect 1662 468 1666 472
rect 30 459 34 463
rect 62 458 66 462
rect 126 458 130 462
rect 150 458 154 462
rect 158 458 162 462
rect 278 458 282 462
rect 286 458 290 462
rect 382 459 386 463
rect 542 458 546 462
rect 574 458 578 462
rect 582 458 586 462
rect 638 458 642 462
rect 662 458 666 462
rect 686 458 690 462
rect 750 458 754 462
rect 838 458 842 462
rect 918 458 922 462
rect 926 458 930 462
rect 982 458 986 462
rect 1014 458 1018 462
rect 1022 458 1026 462
rect 1054 458 1058 462
rect 1126 458 1130 462
rect 1206 458 1210 462
rect 1246 458 1250 462
rect 1278 458 1282 462
rect 1302 458 1306 462
rect 1310 458 1314 462
rect 1334 458 1338 462
rect 1342 458 1346 462
rect 1366 458 1370 462
rect 1486 458 1490 462
rect 1494 458 1498 462
rect 1518 458 1522 462
rect 1542 458 1546 462
rect 1598 458 1602 462
rect 1614 458 1618 462
rect 1670 458 1674 462
rect 1742 458 1746 462
rect 1766 458 1770 462
rect 198 448 202 452
rect 1190 448 1194 452
rect 1262 448 1266 452
rect 1558 448 1562 452
rect 1686 448 1690 452
rect 878 438 882 442
rect 110 418 114 422
rect 1070 418 1074 422
rect 1358 418 1362 422
rect 1510 418 1514 422
rect 1710 418 1714 422
rect 370 403 374 407
rect 377 403 381 407
rect 1386 403 1390 407
rect 1393 403 1397 407
rect 94 388 98 392
rect 174 388 178 392
rect 446 388 450 392
rect 502 388 506 392
rect 550 388 554 392
rect 598 388 602 392
rect 654 388 658 392
rect 718 388 722 392
rect 814 388 818 392
rect 1038 388 1042 392
rect 1206 388 1210 392
rect 1254 388 1258 392
rect 1422 388 1426 392
rect 1462 388 1466 392
rect 1582 388 1586 392
rect 1766 388 1770 392
rect 278 368 282 372
rect 438 368 442 372
rect 798 378 802 382
rect 478 368 482 372
rect 510 368 514 372
rect 558 368 562 372
rect 646 368 650 372
rect 838 368 842 372
rect 1102 368 1106 372
rect 462 358 466 362
rect 542 358 546 362
rect 662 358 666 362
rect 734 358 738 362
rect 910 358 914 362
rect 1222 358 1226 362
rect 1430 358 1434 362
rect 38 348 42 352
rect 110 348 114 352
rect 134 348 138 352
rect 142 348 146 352
rect 150 348 154 352
rect 182 348 186 352
rect 222 348 226 352
rect 286 348 290 352
rect 294 348 298 352
rect 350 348 354 352
rect 358 348 362 352
rect 446 348 450 352
rect 470 348 474 352
rect 494 348 498 352
rect 502 348 506 352
rect 550 348 554 352
rect 574 348 578 352
rect 590 348 594 352
rect 694 348 698 352
rect 726 348 730 352
rect 758 348 762 352
rect 798 348 802 352
rect 806 348 810 352
rect 830 348 834 352
rect 870 348 874 352
rect 886 348 890 352
rect 894 348 898 352
rect 974 347 978 351
rect 1062 348 1066 352
rect 1094 348 1098 352
rect 1142 348 1146 352
rect 1206 348 1210 352
rect 1358 347 1362 351
rect 1462 348 1466 352
rect 1510 348 1514 352
rect 1622 348 1626 352
rect 1638 348 1642 352
rect 1646 348 1650 352
rect 1694 348 1698 352
rect 1710 348 1714 352
rect 1750 348 1754 352
rect 1758 348 1762 352
rect 1782 348 1786 352
rect 102 338 106 342
rect 158 338 162 342
rect 174 338 178 342
rect 526 338 530 342
rect 534 338 538 342
rect 622 338 626 342
rect 646 338 650 342
rect 686 338 690 342
rect 750 338 754 342
rect 774 338 778 342
rect 838 338 842 342
rect 854 338 858 342
rect 958 338 962 342
rect 1086 338 1090 342
rect 1158 338 1162 342
rect 1198 338 1202 342
rect 1238 338 1242 342
rect 1326 338 1330 342
rect 1342 338 1346 342
rect 1470 338 1474 342
rect 1502 338 1506 342
rect 30 328 34 332
rect 214 328 218 332
rect 302 328 306 332
rect 342 328 346 332
rect 422 328 426 332
rect 590 328 594 332
rect 622 328 626 332
rect 678 328 682 332
rect 774 328 778 332
rect 822 328 826 332
rect 942 328 946 332
rect 1046 328 1050 332
rect 1078 328 1082 332
rect 1230 328 1234 332
rect 1590 328 1594 332
rect 374 318 378 322
rect 790 318 794 322
rect 1254 318 1258 322
rect 1270 318 1274 322
rect 1654 318 1658 322
rect 890 303 894 307
rect 897 303 901 307
rect 94 288 98 292
rect 190 288 194 292
rect 214 288 218 292
rect 366 288 370 292
rect 406 288 410 292
rect 454 288 458 292
rect 534 288 538 292
rect 574 288 578 292
rect 654 288 658 292
rect 686 288 690 292
rect 758 288 762 292
rect 798 288 802 292
rect 822 288 826 292
rect 1166 288 1170 292
rect 1254 288 1258 292
rect 1366 288 1370 292
rect 1422 288 1426 292
rect 1454 288 1458 292
rect 1558 288 1562 292
rect 1566 288 1570 292
rect 1694 288 1698 292
rect 1702 288 1706 292
rect 1718 288 1722 292
rect 1774 288 1778 292
rect 30 278 34 282
rect 590 278 594 282
rect 638 278 642 282
rect 678 278 682 282
rect 710 278 714 282
rect 766 278 770 282
rect 814 278 818 282
rect 918 278 922 282
rect 1054 278 1058 282
rect 1238 278 1242 282
rect 1438 278 1442 282
rect 1550 278 1554 282
rect 1598 278 1602 282
rect 1710 278 1714 282
rect 118 268 122 272
rect 174 268 178 272
rect 190 268 194 272
rect 270 268 274 272
rect 286 268 290 272
rect 374 268 378 272
rect 414 268 418 272
rect 446 268 450 272
rect 470 268 474 272
rect 38 258 42 262
rect 62 258 66 262
rect 150 258 154 262
rect 158 258 162 262
rect 166 258 170 262
rect 198 258 202 262
rect 310 258 314 262
rect 334 258 338 262
rect 406 258 410 262
rect 446 258 450 262
rect 494 258 498 262
rect 518 258 522 262
rect 542 258 546 262
rect 558 268 562 272
rect 598 268 602 272
rect 622 268 626 272
rect 702 268 706 272
rect 758 268 762 272
rect 878 268 882 272
rect 950 268 954 272
rect 1038 268 1042 272
rect 1142 268 1146 272
rect 1174 268 1178 272
rect 1222 268 1226 272
rect 1262 268 1266 272
rect 1390 268 1394 272
rect 1582 268 1586 272
rect 1614 268 1618 272
rect 1742 268 1746 272
rect 1798 268 1802 272
rect 750 258 754 262
rect 774 258 778 262
rect 798 258 802 262
rect 886 259 890 263
rect 982 258 986 262
rect 998 258 1002 262
rect 1006 258 1010 262
rect 1118 258 1122 262
rect 1182 258 1186 262
rect 1190 258 1194 262
rect 1302 258 1306 262
rect 1326 258 1330 262
rect 1406 258 1410 262
rect 1494 258 1498 262
rect 1510 258 1514 262
rect 1646 258 1650 262
rect 1734 258 1738 262
rect 1758 258 1762 262
rect 454 248 458 252
rect 502 248 506 252
rect 510 248 514 252
rect 614 248 618 252
rect 646 248 650 252
rect 1158 248 1162 252
rect 1246 248 1250 252
rect 1366 248 1370 252
rect 1414 248 1418 252
rect 1566 248 1570 252
rect 1718 248 1722 252
rect 1782 248 1786 252
rect 422 238 426 242
rect 486 238 490 242
rect 494 238 498 242
rect 598 238 602 242
rect 494 218 498 222
rect 1446 218 1450 222
rect 1590 218 1594 222
rect 370 203 374 207
rect 377 203 381 207
rect 1386 203 1390 207
rect 1393 203 1397 207
rect 126 188 130 192
rect 462 188 466 192
rect 686 188 690 192
rect 782 188 786 192
rect 798 188 802 192
rect 974 188 978 192
rect 1366 188 1370 192
rect 1462 188 1466 192
rect 1622 188 1626 192
rect 1646 188 1650 192
rect 1686 188 1690 192
rect 1734 188 1738 192
rect 142 168 146 172
rect 374 168 378 172
rect 62 158 66 162
rect 678 158 682 162
rect 1102 158 1106 162
rect 1134 158 1138 162
rect 1694 158 1698 162
rect 1710 158 1714 162
rect 1718 158 1722 162
rect 14 148 18 152
rect 38 148 42 152
rect 46 148 50 152
rect 70 148 74 152
rect 102 148 106 152
rect 190 147 194 151
rect 222 148 226 152
rect 230 148 234 152
rect 318 148 322 152
rect 334 148 338 152
rect 398 148 402 152
rect 406 148 410 152
rect 526 147 530 151
rect 574 148 578 152
rect 606 148 610 152
rect 662 148 666 152
rect 670 148 674 152
rect 718 148 722 152
rect 750 148 754 152
rect 862 147 866 151
rect 958 148 962 152
rect 966 148 970 152
rect 1006 148 1010 152
rect 1038 147 1042 151
rect 1118 148 1122 152
rect 1126 148 1130 152
rect 1150 148 1154 152
rect 1158 148 1162 152
rect 1182 148 1186 152
rect 1198 148 1202 152
rect 1214 148 1218 152
rect 1222 148 1226 152
rect 1246 148 1250 152
rect 1294 148 1298 152
rect 1406 148 1410 152
rect 1430 148 1434 152
rect 1446 148 1450 152
rect 1470 148 1474 152
rect 1478 148 1482 152
rect 1486 148 1490 152
rect 1494 148 1498 152
rect 1526 148 1530 152
rect 1558 147 1562 151
rect 1582 148 1586 152
rect 1630 148 1634 152
rect 1638 148 1642 152
rect 1662 148 1666 152
rect 1758 148 1762 152
rect 1782 148 1786 152
rect 1790 148 1794 152
rect 78 138 82 142
rect 182 138 186 142
rect 294 138 298 142
rect 446 138 450 142
rect 598 138 602 142
rect 630 138 634 142
rect 694 138 698 142
rect 742 138 746 142
rect 790 138 794 142
rect 830 138 834 142
rect 878 138 882 142
rect 926 138 930 142
rect 1270 138 1274 142
rect 1382 138 1386 142
rect 1518 138 1522 142
rect 1542 138 1546 142
rect 1678 138 1682 142
rect 62 128 66 132
rect 118 128 122 132
rect 158 128 162 132
rect 278 128 282 132
rect 414 128 418 132
rect 494 128 498 132
rect 526 128 530 132
rect 558 128 562 132
rect 590 128 594 132
rect 614 128 618 132
rect 910 128 914 132
rect 1070 128 1074 132
rect 1134 128 1138 132
rect 1198 128 1202 132
rect 1710 128 1714 132
rect 1718 128 1722 132
rect 1742 128 1746 132
rect 30 118 34 122
rect 86 118 90 122
rect 246 118 250 122
rect 734 118 738 122
rect 1166 118 1170 122
rect 1230 118 1234 122
rect 1766 118 1770 122
rect 890 103 894 107
rect 897 103 901 107
rect 94 88 98 92
rect 190 88 194 92
rect 214 88 218 92
rect 342 88 346 92
rect 454 88 458 92
rect 606 88 610 92
rect 638 88 642 92
rect 654 88 658 92
rect 838 88 842 92
rect 950 88 954 92
rect 966 88 970 92
rect 1070 88 1074 92
rect 1174 88 1178 92
rect 1230 88 1234 92
rect 1366 88 1370 92
rect 1598 88 1602 92
rect 1694 88 1698 92
rect 1790 88 1794 92
rect 46 68 50 72
rect 110 68 114 72
rect 142 68 146 72
rect 206 68 210 72
rect 230 78 234 82
rect 494 78 498 82
rect 1222 78 1226 82
rect 1254 78 1258 82
rect 1382 78 1386 82
rect 294 68 298 72
rect 374 68 378 72
rect 502 68 506 72
rect 526 68 530 72
rect 646 68 650 72
rect 782 68 786 72
rect 862 68 866 72
rect 958 68 962 72
rect 1046 68 1050 72
rect 1078 68 1082 72
rect 1118 68 1122 72
rect 1214 68 1218 72
rect 1270 68 1274 72
rect 1358 68 1362 72
rect 1398 68 1402 72
rect 1502 68 1506 72
rect 1542 68 1546 72
rect 1614 68 1618 72
rect 1710 68 1714 72
rect 30 59 34 63
rect 126 59 130 63
rect 198 58 202 62
rect 246 58 250 62
rect 278 59 282 63
rect 414 58 418 62
rect 478 58 482 62
rect 510 58 514 62
rect 550 58 554 62
rect 718 59 722 63
rect 782 58 786 62
rect 894 58 898 62
rect 902 58 906 62
rect 926 58 930 62
rect 1030 59 1034 63
rect 1126 58 1130 62
rect 1214 58 1218 62
rect 1294 58 1298 62
rect 1446 58 1450 62
rect 1462 58 1466 62
rect 1470 58 1474 62
rect 1494 58 1498 62
rect 1534 59 1538 63
rect 1638 58 1642 62
rect 1726 59 1730 63
rect 1374 48 1378 52
rect 1062 38 1066 42
rect 370 3 374 7
rect 377 3 381 7
rect 1386 3 1390 7
rect 1393 3 1397 7
<< metal2 >>
rect 598 1728 602 1732
rect 718 1728 722 1732
rect 830 1728 834 1732
rect 870 1728 874 1732
rect 1302 1728 1306 1732
rect 154 1688 158 1691
rect 522 1688 526 1691
rect 14 1682 17 1688
rect 62 1662 65 1668
rect 38 1652 41 1658
rect 54 1552 57 1658
rect 94 1652 97 1659
rect 126 1612 129 1658
rect 62 1552 65 1608
rect 38 1542 41 1548
rect 62 1462 65 1548
rect 102 1532 105 1568
rect 150 1552 153 1618
rect 206 1592 209 1658
rect 222 1612 225 1658
rect 186 1558 190 1561
rect 202 1548 206 1551
rect 122 1538 126 1541
rect 106 1528 110 1531
rect 94 1482 97 1488
rect 106 1478 110 1481
rect 138 1468 142 1471
rect 118 1462 121 1468
rect 126 1462 129 1468
rect 150 1462 153 1548
rect 158 1542 161 1548
rect 190 1542 193 1548
rect 166 1532 169 1538
rect 158 1472 161 1478
rect 42 1458 46 1461
rect 62 1352 65 1458
rect 150 1362 153 1458
rect 174 1442 177 1448
rect 182 1442 185 1518
rect 202 1478 206 1481
rect 222 1462 225 1548
rect 254 1542 257 1618
rect 262 1592 265 1618
rect 286 1592 289 1608
rect 266 1558 270 1561
rect 254 1462 257 1468
rect 190 1452 193 1458
rect 194 1368 198 1371
rect 206 1352 209 1358
rect 138 1348 142 1351
rect 30 1292 33 1347
rect 62 1342 65 1348
rect 110 1342 113 1348
rect 46 1262 49 1318
rect 94 1312 97 1318
rect 62 1282 65 1308
rect 158 1282 161 1338
rect 198 1322 201 1348
rect 122 1278 126 1281
rect 110 1262 113 1268
rect 18 1258 22 1261
rect 58 1258 62 1261
rect 38 1252 41 1258
rect 26 1168 30 1171
rect 38 1152 41 1158
rect 46 1152 49 1238
rect 70 1192 73 1258
rect 78 1162 81 1258
rect 18 1148 22 1151
rect 58 1148 62 1151
rect 94 1151 97 1168
rect 38 1052 41 1058
rect 34 948 38 951
rect 30 882 33 928
rect 34 858 38 861
rect 34 748 38 751
rect 6 652 9 668
rect 18 548 22 551
rect 30 542 33 618
rect 38 552 41 728
rect 46 662 49 1148
rect 62 1132 65 1138
rect 62 1062 65 1088
rect 102 1062 105 1248
rect 126 1152 129 1268
rect 158 1252 161 1259
rect 214 1252 217 1458
rect 222 1362 225 1458
rect 270 1382 273 1518
rect 254 1362 257 1368
rect 226 1348 230 1351
rect 222 1282 225 1288
rect 230 1252 233 1308
rect 238 1262 241 1348
rect 254 1332 257 1358
rect 262 1321 265 1368
rect 278 1362 281 1418
rect 286 1392 289 1448
rect 318 1362 321 1688
rect 430 1682 433 1688
rect 342 1672 345 1678
rect 598 1672 601 1728
rect 718 1682 721 1728
rect 830 1682 833 1728
rect 870 1682 873 1728
rect 888 1703 890 1707
rect 894 1703 897 1707
rect 901 1703 904 1707
rect 1254 1682 1257 1688
rect 702 1672 705 1678
rect 814 1672 817 1678
rect 854 1672 857 1678
rect 414 1662 417 1668
rect 326 1582 329 1659
rect 370 1658 374 1661
rect 382 1642 385 1658
rect 342 1542 345 1628
rect 368 1603 370 1607
rect 374 1603 377 1607
rect 381 1603 384 1607
rect 422 1552 425 1668
rect 494 1662 497 1668
rect 462 1652 465 1659
rect 538 1658 542 1661
rect 598 1632 601 1668
rect 614 1662 617 1668
rect 638 1592 641 1658
rect 538 1578 542 1581
rect 358 1472 361 1538
rect 398 1522 401 1548
rect 422 1502 425 1548
rect 478 1542 481 1548
rect 498 1538 502 1541
rect 446 1518 454 1521
rect 402 1468 406 1471
rect 422 1462 425 1468
rect 330 1458 334 1461
rect 390 1432 393 1458
rect 418 1448 422 1451
rect 368 1403 370 1407
rect 374 1403 377 1407
rect 381 1403 384 1407
rect 366 1372 369 1378
rect 338 1368 342 1371
rect 306 1358 310 1361
rect 274 1348 278 1351
rect 294 1342 297 1358
rect 330 1348 334 1351
rect 310 1342 313 1348
rect 358 1342 361 1348
rect 386 1328 390 1331
rect 254 1318 265 1321
rect 158 1152 161 1168
rect 166 1152 169 1158
rect 126 1092 129 1148
rect 158 1132 161 1148
rect 198 1142 201 1148
rect 178 1138 182 1141
rect 114 1068 118 1071
rect 134 1062 137 1068
rect 122 1058 126 1061
rect 94 1022 97 1028
rect 94 972 97 978
rect 102 942 105 1058
rect 134 982 137 1058
rect 150 1022 153 1078
rect 166 1072 169 1088
rect 182 1063 185 1118
rect 198 1072 201 1138
rect 206 1082 209 1248
rect 254 1242 257 1318
rect 354 1288 358 1291
rect 250 1238 254 1241
rect 254 1182 257 1218
rect 270 1152 273 1268
rect 294 1262 297 1268
rect 318 1152 321 1158
rect 350 1152 353 1278
rect 374 1262 377 1318
rect 390 1272 393 1278
rect 386 1258 390 1261
rect 374 1222 377 1258
rect 368 1203 370 1207
rect 374 1203 377 1207
rect 381 1203 384 1207
rect 398 1192 401 1228
rect 254 1132 257 1148
rect 350 1142 353 1148
rect 366 1142 369 1148
rect 214 1082 217 1128
rect 150 962 153 1018
rect 158 952 161 988
rect 166 952 169 958
rect 146 948 150 951
rect 118 942 121 948
rect 98 888 102 891
rect 106 878 110 881
rect 118 872 121 898
rect 102 862 105 868
rect 126 862 129 948
rect 150 882 153 888
rect 174 882 177 938
rect 182 892 185 978
rect 198 952 201 978
rect 210 948 214 951
rect 206 932 209 938
rect 138 878 142 881
rect 174 862 177 868
rect 62 752 65 858
rect 126 811 129 858
rect 178 848 182 851
rect 118 808 129 811
rect 62 722 65 748
rect 94 722 97 738
rect 118 732 121 808
rect 126 772 129 778
rect 102 702 105 718
rect 54 662 57 668
rect 78 662 81 668
rect 86 662 89 698
rect 110 692 113 728
rect 98 688 102 691
rect 46 572 49 658
rect 46 552 49 568
rect 70 552 73 558
rect 58 548 62 551
rect 30 463 33 518
rect 38 362 41 548
rect 94 542 97 588
rect 134 562 137 758
rect 158 742 161 748
rect 142 732 145 738
rect 146 728 150 731
rect 158 672 161 718
rect 182 692 185 818
rect 190 762 193 918
rect 214 902 217 948
rect 222 922 225 928
rect 206 872 209 878
rect 218 868 222 871
rect 198 862 201 868
rect 230 852 233 1118
rect 246 1092 249 1128
rect 310 1112 313 1118
rect 326 1111 329 1138
rect 338 1128 342 1131
rect 366 1122 369 1128
rect 318 1108 329 1111
rect 278 1072 281 1078
rect 302 1072 305 1088
rect 262 1051 265 1068
rect 262 1048 273 1051
rect 238 952 241 958
rect 246 942 249 948
rect 254 942 257 948
rect 246 932 249 938
rect 258 918 262 921
rect 254 882 257 888
rect 270 882 273 1048
rect 278 1032 281 1038
rect 286 1021 289 1058
rect 278 1018 289 1021
rect 258 858 262 861
rect 278 852 281 1018
rect 302 952 305 958
rect 286 862 289 888
rect 294 872 297 948
rect 274 848 278 851
rect 214 792 217 838
rect 222 782 225 818
rect 198 752 201 778
rect 230 772 233 848
rect 242 838 246 841
rect 254 792 257 838
rect 262 792 265 848
rect 302 842 305 878
rect 278 822 281 828
rect 242 768 246 771
rect 218 758 222 761
rect 230 752 233 758
rect 298 748 302 751
rect 310 751 313 938
rect 318 932 321 1108
rect 386 1088 390 1091
rect 398 1062 401 1178
rect 406 1162 409 1388
rect 326 1052 329 1058
rect 326 861 329 1018
rect 368 1003 370 1007
rect 374 1003 377 1007
rect 381 1003 384 1007
rect 378 968 382 971
rect 358 962 361 968
rect 366 952 369 958
rect 322 858 329 861
rect 338 859 345 861
rect 338 858 342 859
rect 350 852 353 858
rect 366 842 369 918
rect 374 862 377 908
rect 390 842 393 868
rect 350 792 353 838
rect 398 822 401 1058
rect 406 1042 409 1158
rect 414 1152 417 1218
rect 422 1152 425 1428
rect 430 1342 433 1498
rect 438 1482 441 1488
rect 446 1472 449 1518
rect 478 1472 481 1538
rect 498 1518 502 1521
rect 510 1512 513 1548
rect 518 1532 521 1548
rect 518 1502 521 1528
rect 494 1482 497 1498
rect 462 1442 465 1448
rect 430 1332 433 1338
rect 430 1282 433 1288
rect 438 1272 441 1348
rect 454 1312 457 1418
rect 478 1352 481 1468
rect 494 1463 497 1468
rect 526 1462 529 1548
rect 574 1542 577 1588
rect 602 1558 606 1561
rect 678 1552 681 1638
rect 742 1632 745 1668
rect 882 1658 886 1661
rect 806 1652 809 1658
rect 878 1642 881 1658
rect 918 1652 921 1668
rect 1046 1662 1049 1668
rect 1018 1658 1022 1661
rect 1114 1658 1118 1661
rect 942 1652 945 1658
rect 1006 1642 1009 1658
rect 1002 1618 1009 1621
rect 694 1612 697 1618
rect 726 1582 729 1618
rect 702 1552 705 1558
rect 602 1548 606 1551
rect 562 1488 566 1491
rect 542 1352 545 1458
rect 574 1392 577 1458
rect 590 1442 593 1518
rect 614 1512 617 1548
rect 726 1542 729 1548
rect 766 1542 769 1548
rect 790 1542 793 1548
rect 806 1542 809 1558
rect 826 1547 830 1550
rect 642 1538 646 1541
rect 778 1538 785 1541
rect 598 1472 601 1488
rect 626 1478 630 1481
rect 634 1468 638 1471
rect 646 1462 649 1478
rect 666 1468 670 1471
rect 610 1448 614 1451
rect 562 1368 566 1371
rect 582 1362 585 1418
rect 606 1362 609 1418
rect 654 1382 657 1448
rect 618 1368 622 1371
rect 654 1362 657 1378
rect 662 1362 665 1368
rect 594 1358 598 1361
rect 498 1348 502 1351
rect 534 1342 537 1348
rect 522 1338 526 1341
rect 490 1318 494 1321
rect 446 1262 449 1308
rect 494 1282 497 1318
rect 510 1302 513 1328
rect 526 1282 529 1328
rect 534 1282 537 1338
rect 454 1272 457 1278
rect 438 1252 441 1258
rect 434 1168 438 1171
rect 446 1162 449 1258
rect 502 1151 505 1168
rect 414 1072 417 1148
rect 422 1142 425 1148
rect 422 1132 425 1138
rect 470 1132 473 1148
rect 510 1142 513 1268
rect 534 1262 537 1268
rect 542 1262 545 1348
rect 518 1131 521 1218
rect 550 1162 553 1358
rect 558 1342 561 1348
rect 582 1322 585 1338
rect 614 1332 617 1348
rect 678 1342 681 1488
rect 686 1432 689 1528
rect 734 1512 737 1528
rect 686 1342 689 1408
rect 702 1362 705 1388
rect 718 1352 721 1358
rect 734 1352 737 1508
rect 750 1482 753 1538
rect 782 1462 785 1538
rect 790 1492 793 1528
rect 750 1392 753 1459
rect 774 1362 777 1388
rect 758 1352 761 1358
rect 782 1352 785 1458
rect 798 1452 801 1478
rect 806 1462 809 1498
rect 838 1462 841 1618
rect 930 1588 934 1591
rect 906 1548 910 1551
rect 918 1532 921 1548
rect 1006 1532 1009 1618
rect 1070 1572 1073 1618
rect 1126 1572 1129 1668
rect 1174 1592 1177 1618
rect 1146 1568 1150 1571
rect 1014 1562 1017 1568
rect 1018 1548 1022 1551
rect 966 1522 969 1528
rect 974 1522 977 1528
rect 878 1518 886 1521
rect 846 1462 849 1468
rect 818 1458 822 1461
rect 878 1452 881 1518
rect 888 1503 890 1507
rect 894 1503 897 1507
rect 901 1503 904 1507
rect 930 1468 934 1471
rect 938 1458 942 1461
rect 982 1452 985 1498
rect 990 1482 993 1488
rect 998 1462 1001 1468
rect 1006 1462 1009 1528
rect 1022 1502 1025 1548
rect 1030 1542 1033 1548
rect 1014 1492 1017 1498
rect 1014 1472 1017 1478
rect 726 1342 729 1348
rect 590 1292 593 1298
rect 598 1262 601 1318
rect 606 1272 609 1278
rect 614 1272 617 1328
rect 610 1258 614 1261
rect 622 1252 625 1318
rect 638 1302 641 1338
rect 678 1332 681 1338
rect 714 1328 718 1331
rect 734 1322 737 1348
rect 790 1342 793 1418
rect 798 1362 801 1378
rect 806 1351 809 1428
rect 798 1348 809 1351
rect 630 1252 633 1288
rect 638 1262 641 1268
rect 646 1252 649 1318
rect 670 1302 673 1318
rect 702 1311 705 1318
rect 702 1308 713 1311
rect 678 1262 681 1268
rect 658 1258 662 1261
rect 686 1252 689 1268
rect 702 1262 705 1298
rect 710 1242 713 1308
rect 758 1282 761 1288
rect 730 1258 734 1261
rect 722 1248 726 1251
rect 742 1242 745 1248
rect 642 1238 646 1241
rect 666 1238 670 1241
rect 606 1232 609 1238
rect 718 1172 721 1218
rect 566 1152 569 1168
rect 726 1152 729 1228
rect 766 1222 769 1268
rect 774 1252 777 1318
rect 798 1292 801 1348
rect 814 1342 817 1448
rect 882 1418 886 1421
rect 922 1358 926 1361
rect 850 1348 854 1351
rect 874 1348 878 1351
rect 826 1328 830 1331
rect 786 1258 790 1261
rect 714 1148 718 1151
rect 510 1128 521 1131
rect 462 1082 465 1088
rect 462 1072 465 1078
rect 470 1072 473 1118
rect 510 1092 513 1128
rect 542 1092 545 1098
rect 574 1082 577 1118
rect 630 1112 633 1148
rect 654 1132 657 1138
rect 598 1092 601 1108
rect 670 1091 673 1128
rect 670 1088 678 1091
rect 578 1078 582 1081
rect 550 1072 553 1078
rect 530 1068 534 1071
rect 558 1062 561 1078
rect 670 1072 673 1088
rect 418 1058 422 1061
rect 494 1058 502 1061
rect 474 1048 478 1051
rect 430 1042 433 1048
rect 486 1032 489 1048
rect 494 1032 497 1058
rect 514 1048 518 1051
rect 506 1038 510 1041
rect 454 992 457 998
rect 478 992 481 1008
rect 510 992 513 1028
rect 406 942 409 978
rect 418 948 422 951
rect 446 942 449 968
rect 462 962 465 978
rect 474 958 478 961
rect 474 948 478 951
rect 454 941 457 948
rect 454 938 462 941
rect 406 922 409 938
rect 422 892 425 938
rect 430 922 433 928
rect 454 892 457 928
rect 474 888 478 891
rect 434 868 438 871
rect 446 862 449 868
rect 406 852 409 858
rect 368 803 370 807
rect 374 803 377 807
rect 381 803 384 807
rect 390 802 393 818
rect 310 748 318 751
rect 190 741 193 748
rect 190 738 201 741
rect 198 672 201 738
rect 206 732 209 738
rect 238 692 241 748
rect 278 682 281 688
rect 286 682 289 688
rect 266 678 270 681
rect 254 672 257 678
rect 266 668 270 671
rect 146 658 150 661
rect 158 551 161 668
rect 198 662 201 668
rect 222 662 225 668
rect 238 662 241 668
rect 190 652 193 658
rect 198 652 201 658
rect 62 462 65 528
rect 78 492 81 538
rect 86 452 89 518
rect 94 492 97 498
rect 102 482 105 548
rect 158 548 166 551
rect 134 492 137 547
rect 166 532 169 548
rect 174 482 177 508
rect 190 492 193 638
rect 214 592 217 658
rect 238 592 241 648
rect 206 562 209 588
rect 226 568 230 571
rect 278 562 281 568
rect 222 542 225 548
rect 246 542 249 558
rect 286 552 289 678
rect 318 662 321 748
rect 374 742 377 748
rect 390 692 393 778
rect 382 662 385 668
rect 330 658 334 661
rect 198 512 201 518
rect 102 391 105 478
rect 166 472 169 478
rect 126 462 129 468
rect 162 458 166 461
rect 150 442 153 458
rect 98 388 105 391
rect 110 352 113 418
rect 134 352 137 358
rect 142 352 145 398
rect 174 392 177 468
rect 194 448 198 451
rect 206 432 209 518
rect 214 492 217 528
rect 206 402 209 428
rect 182 352 185 358
rect 42 348 46 351
rect 102 342 105 348
rect 30 282 33 328
rect 94 292 97 298
rect 62 262 65 288
rect 118 262 121 268
rect 42 258 46 261
rect 14 152 17 158
rect 38 152 41 248
rect 126 192 129 268
rect 134 252 137 348
rect 150 272 153 348
rect 222 342 225 348
rect 158 282 161 338
rect 174 302 177 338
rect 190 292 193 318
rect 214 292 217 328
rect 174 272 177 278
rect 158 262 161 268
rect 150 252 153 258
rect 46 152 49 168
rect 58 158 62 161
rect 66 148 70 151
rect 78 142 81 148
rect 30 63 33 118
rect 62 92 65 128
rect 50 68 54 71
rect 86 62 89 118
rect 94 102 97 178
rect 106 148 110 151
rect 122 128 126 131
rect 94 92 97 98
rect 110 72 113 78
rect 142 72 145 168
rect 166 132 169 258
rect 182 142 185 288
rect 230 271 233 458
rect 254 442 257 548
rect 262 542 265 548
rect 222 268 233 271
rect 190 182 193 268
rect 202 258 206 261
rect 222 172 225 268
rect 222 152 225 168
rect 230 152 233 248
rect 158 82 161 128
rect 166 102 169 128
rect 190 122 193 147
rect 190 92 193 98
rect 126 63 129 68
rect 198 62 201 108
rect 206 72 209 148
rect 214 92 217 118
rect 230 112 233 148
rect 226 78 230 81
rect 246 72 249 118
rect 206 62 209 68
rect 262 62 265 538
rect 302 532 305 548
rect 318 542 321 658
rect 406 621 409 848
rect 430 752 433 818
rect 438 782 441 858
rect 462 842 465 848
rect 446 792 449 838
rect 454 752 457 758
rect 422 711 425 748
rect 438 722 441 738
rect 422 708 433 711
rect 422 662 425 668
rect 430 662 433 708
rect 470 672 473 738
rect 486 692 489 968
rect 502 962 505 978
rect 502 762 505 958
rect 518 902 521 938
rect 518 892 521 898
rect 526 852 529 1058
rect 566 1052 569 1058
rect 574 952 577 1068
rect 606 1052 609 1068
rect 654 1062 657 1068
rect 634 1058 638 1061
rect 614 1012 617 1058
rect 650 1048 654 1051
rect 622 972 625 1048
rect 694 1042 697 1128
rect 710 1061 713 1118
rect 710 1058 718 1061
rect 642 1038 646 1041
rect 630 1022 633 1028
rect 678 992 681 1018
rect 646 952 649 968
rect 626 948 630 951
rect 702 942 705 948
rect 562 938 566 941
rect 578 928 582 931
rect 598 922 601 938
rect 534 863 537 888
rect 550 872 553 918
rect 566 882 569 918
rect 586 888 590 891
rect 598 882 601 898
rect 646 892 649 908
rect 622 872 625 888
rect 702 882 705 898
rect 726 881 729 1148
rect 734 1002 737 1138
rect 742 1132 745 1168
rect 750 1152 753 1218
rect 806 1181 809 1318
rect 838 1312 841 1338
rect 878 1322 881 1338
rect 890 1318 894 1321
rect 814 1192 817 1308
rect 888 1303 890 1307
rect 894 1303 897 1307
rect 901 1303 904 1307
rect 854 1272 857 1278
rect 862 1262 865 1268
rect 806 1178 817 1181
rect 758 1132 761 1148
rect 782 1082 785 1148
rect 778 1068 782 1071
rect 758 1041 761 1068
rect 758 1038 769 1041
rect 766 972 769 1038
rect 790 1032 793 1118
rect 806 1102 809 1168
rect 814 1162 817 1178
rect 830 1162 833 1168
rect 926 1162 929 1348
rect 934 1342 937 1418
rect 958 1352 961 1388
rect 954 1338 958 1341
rect 1014 1332 1017 1468
rect 1038 1392 1041 1518
rect 1046 1472 1049 1518
rect 1054 1472 1057 1568
rect 1094 1552 1097 1558
rect 1186 1548 1190 1551
rect 1086 1482 1089 1488
rect 1070 1472 1073 1478
rect 1086 1462 1089 1478
rect 1102 1472 1105 1528
rect 1118 1492 1121 1548
rect 1254 1542 1257 1648
rect 1134 1492 1137 1518
rect 1142 1462 1145 1538
rect 1150 1462 1153 1508
rect 1158 1462 1161 1498
rect 1190 1472 1193 1538
rect 1270 1532 1273 1668
rect 1302 1662 1305 1728
rect 1550 1692 1553 1698
rect 1438 1682 1441 1688
rect 1766 1682 1769 1688
rect 1566 1672 1569 1678
rect 1422 1662 1425 1668
rect 1322 1658 1326 1661
rect 1366 1652 1369 1658
rect 1318 1622 1321 1648
rect 1278 1552 1281 1578
rect 1302 1552 1305 1578
rect 1234 1528 1238 1531
rect 1130 1458 1134 1461
rect 1030 1351 1033 1368
rect 1046 1352 1049 1458
rect 1070 1382 1073 1418
rect 1078 1352 1081 1358
rect 1142 1352 1145 1458
rect 1150 1382 1153 1458
rect 1174 1442 1177 1448
rect 1066 1348 1070 1351
rect 1026 1338 1030 1341
rect 926 1152 929 1158
rect 850 1148 854 1151
rect 814 1122 817 1148
rect 862 1142 865 1148
rect 910 1142 913 1148
rect 934 1142 937 1238
rect 942 1172 945 1318
rect 966 1282 969 1318
rect 1038 1292 1041 1298
rect 1070 1292 1073 1338
rect 1086 1332 1089 1338
rect 1102 1332 1105 1348
rect 1102 1302 1105 1328
rect 1078 1292 1081 1298
rect 1066 1278 1070 1281
rect 954 1268 958 1271
rect 966 1212 969 1278
rect 1018 1268 1022 1271
rect 998 1262 1001 1268
rect 1030 1262 1033 1268
rect 1134 1262 1137 1318
rect 1150 1312 1153 1348
rect 1158 1342 1161 1348
rect 1190 1342 1193 1468
rect 1246 1462 1249 1468
rect 1270 1452 1273 1458
rect 1210 1418 1214 1421
rect 1278 1392 1281 1548
rect 1286 1542 1289 1548
rect 1294 1512 1297 1548
rect 1334 1542 1337 1548
rect 1350 1522 1353 1528
rect 1358 1511 1361 1648
rect 1390 1631 1393 1650
rect 1384 1603 1386 1607
rect 1390 1603 1393 1607
rect 1397 1603 1400 1607
rect 1398 1551 1401 1558
rect 1478 1552 1481 1658
rect 1466 1538 1470 1541
rect 1350 1508 1361 1511
rect 1310 1472 1313 1478
rect 1342 1462 1345 1468
rect 1350 1462 1353 1508
rect 1398 1482 1401 1528
rect 1314 1458 1318 1461
rect 1362 1458 1366 1461
rect 1278 1352 1281 1388
rect 1318 1361 1321 1458
rect 1326 1452 1329 1458
rect 1326 1361 1329 1368
rect 1318 1358 1329 1361
rect 1326 1352 1329 1358
rect 1342 1352 1345 1358
rect 1266 1348 1270 1351
rect 1306 1348 1310 1351
rect 1198 1342 1201 1348
rect 1282 1338 1286 1341
rect 1190 1332 1193 1338
rect 1170 1288 1174 1291
rect 1238 1282 1241 1328
rect 1270 1282 1273 1288
rect 1158 1272 1161 1278
rect 1206 1272 1209 1278
rect 1274 1268 1278 1271
rect 1238 1263 1241 1268
rect 1058 1258 1062 1261
rect 1294 1262 1297 1308
rect 1310 1302 1313 1348
rect 1318 1332 1321 1348
rect 1350 1332 1353 1458
rect 1384 1403 1386 1407
rect 1390 1403 1393 1407
rect 1397 1403 1400 1407
rect 1362 1348 1369 1351
rect 1306 1278 1310 1281
rect 1366 1272 1369 1348
rect 1354 1268 1358 1271
rect 1318 1262 1321 1268
rect 958 1182 961 1188
rect 958 1142 961 1168
rect 966 1152 969 1168
rect 974 1162 977 1178
rect 850 1138 857 1141
rect 830 1132 833 1138
rect 854 1092 857 1138
rect 930 1128 934 1131
rect 878 1092 881 1118
rect 888 1103 890 1107
rect 894 1103 897 1107
rect 901 1103 904 1107
rect 822 1072 825 1078
rect 734 952 737 958
rect 734 892 737 938
rect 742 922 745 948
rect 750 902 753 918
rect 726 878 737 881
rect 694 872 697 878
rect 682 868 686 871
rect 498 748 502 751
rect 518 682 521 778
rect 534 691 537 798
rect 550 762 553 868
rect 566 862 569 868
rect 574 862 577 868
rect 662 862 665 868
rect 702 862 705 878
rect 618 858 622 861
rect 566 832 569 858
rect 558 762 561 768
rect 574 742 577 768
rect 614 752 617 758
rect 546 718 550 721
rect 558 702 561 718
rect 534 688 545 691
rect 486 672 489 678
rect 506 668 510 671
rect 454 663 457 668
rect 534 662 537 678
rect 542 672 545 688
rect 550 672 553 678
rect 490 658 494 661
rect 566 642 569 658
rect 430 628 438 631
rect 406 618 417 621
rect 368 603 370 607
rect 374 603 377 607
rect 381 603 384 607
rect 334 551 337 558
rect 406 552 409 568
rect 318 532 321 538
rect 350 482 353 488
rect 270 472 273 478
rect 366 472 369 538
rect 414 502 417 618
rect 430 542 433 628
rect 478 592 481 628
rect 526 592 529 598
rect 446 572 449 578
rect 466 568 470 571
rect 498 558 502 561
rect 474 548 478 551
rect 270 272 273 468
rect 278 462 281 468
rect 318 462 321 468
rect 382 463 385 468
rect 286 422 289 458
rect 282 368 286 371
rect 286 352 289 358
rect 294 332 297 348
rect 302 332 305 338
rect 342 332 345 368
rect 350 352 353 358
rect 358 352 361 438
rect 368 403 370 407
rect 374 403 377 407
rect 381 403 384 407
rect 366 292 369 328
rect 374 292 377 318
rect 406 292 409 358
rect 286 272 289 288
rect 310 262 313 288
rect 414 281 417 498
rect 422 332 425 338
rect 406 278 417 281
rect 430 282 433 538
rect 446 512 449 538
rect 454 502 457 548
rect 486 532 489 558
rect 558 552 561 558
rect 566 552 569 568
rect 494 542 497 548
rect 518 542 521 548
rect 526 538 534 541
rect 442 488 446 491
rect 454 472 457 478
rect 454 412 457 468
rect 446 392 449 398
rect 502 392 505 528
rect 510 492 513 528
rect 526 482 529 538
rect 542 532 545 548
rect 534 492 537 498
rect 550 482 553 518
rect 558 492 561 518
rect 526 472 529 478
rect 534 458 542 461
rect 482 368 486 371
rect 438 322 441 368
rect 462 362 465 368
rect 450 348 457 351
rect 454 292 457 348
rect 470 342 473 348
rect 494 332 497 348
rect 502 342 505 348
rect 334 152 337 258
rect 374 222 377 268
rect 406 262 409 278
rect 430 272 433 278
rect 450 268 454 271
rect 318 142 321 148
rect 278 92 281 128
rect 294 72 297 138
rect 342 92 345 218
rect 368 203 370 207
rect 374 203 377 207
rect 381 203 384 207
rect 414 192 417 268
rect 422 242 425 248
rect 374 172 377 188
rect 374 132 377 168
rect 394 148 398 151
rect 410 148 414 151
rect 446 151 449 258
rect 458 248 462 251
rect 470 191 473 268
rect 502 261 505 338
rect 498 258 505 261
rect 510 262 513 368
rect 534 342 537 458
rect 550 392 553 468
rect 554 368 558 371
rect 542 362 545 368
rect 550 352 553 358
rect 526 332 529 338
rect 534 332 537 338
rect 534 292 537 318
rect 550 262 553 288
rect 558 262 561 268
rect 546 258 550 261
rect 486 242 489 258
rect 494 232 497 238
rect 502 232 505 248
rect 510 222 513 248
rect 518 222 521 258
rect 498 218 502 221
rect 466 188 473 191
rect 446 148 457 151
rect 414 132 417 138
rect 446 132 449 138
rect 454 92 457 148
rect 566 151 569 468
rect 574 462 577 708
rect 598 682 601 718
rect 622 672 625 858
rect 642 848 646 851
rect 650 838 654 841
rect 662 822 665 858
rect 678 852 681 858
rect 694 842 697 848
rect 718 822 721 858
rect 630 782 633 818
rect 630 732 633 748
rect 638 692 641 748
rect 646 702 649 728
rect 642 668 646 671
rect 622 662 625 668
rect 662 662 665 758
rect 694 752 697 818
rect 726 752 729 798
rect 734 782 737 878
rect 742 822 745 868
rect 758 862 761 918
rect 798 872 801 1058
rect 822 991 825 1058
rect 830 1022 833 1068
rect 862 1002 865 1068
rect 814 988 825 991
rect 870 991 873 1058
rect 866 988 873 991
rect 814 972 817 988
rect 878 982 881 1048
rect 910 992 913 1068
rect 806 942 809 948
rect 770 858 774 861
rect 750 831 753 858
rect 750 828 761 831
rect 758 812 761 828
rect 742 782 745 788
rect 734 772 737 778
rect 766 772 769 838
rect 734 752 737 768
rect 754 748 758 751
rect 678 732 681 738
rect 694 692 697 748
rect 702 732 705 738
rect 766 701 769 748
rect 774 712 777 858
rect 782 792 785 818
rect 790 792 793 858
rect 806 842 809 848
rect 814 821 817 968
rect 830 932 833 938
rect 842 888 846 891
rect 830 872 833 888
rect 854 882 857 918
rect 888 903 890 907
rect 894 903 897 907
rect 901 903 904 907
rect 910 892 913 948
rect 806 818 817 821
rect 806 752 809 818
rect 822 752 825 868
rect 830 862 833 868
rect 846 852 849 868
rect 918 862 921 948
rect 926 942 929 1018
rect 782 722 785 738
rect 766 698 777 701
rect 670 682 673 688
rect 726 682 729 698
rect 690 668 697 671
rect 678 662 681 668
rect 598 652 601 658
rect 582 472 585 558
rect 598 482 601 488
rect 606 472 609 638
rect 622 562 625 658
rect 666 588 670 591
rect 614 532 617 538
rect 614 482 617 528
rect 622 522 625 548
rect 646 492 649 518
rect 650 468 654 471
rect 662 462 665 548
rect 682 538 686 541
rect 694 532 697 668
rect 738 658 742 661
rect 718 592 721 618
rect 774 602 777 698
rect 794 688 798 691
rect 734 552 737 558
rect 702 542 705 548
rect 674 528 678 531
rect 730 528 734 531
rect 686 492 689 528
rect 634 458 638 461
rect 574 442 577 458
rect 582 431 585 458
rect 574 428 585 431
rect 574 352 577 428
rect 598 392 601 458
rect 654 382 657 388
rect 670 372 673 468
rect 686 462 689 468
rect 646 362 649 368
rect 658 358 662 361
rect 586 348 590 351
rect 574 292 577 348
rect 626 338 630 341
rect 642 338 646 341
rect 594 328 598 331
rect 590 282 593 298
rect 622 282 625 328
rect 630 302 633 338
rect 678 332 681 358
rect 694 352 697 528
rect 702 362 705 478
rect 718 472 721 478
rect 718 392 721 448
rect 686 342 689 348
rect 694 342 697 348
rect 598 272 601 278
rect 618 268 622 271
rect 598 262 601 268
rect 630 262 633 298
rect 638 282 641 318
rect 654 292 657 298
rect 686 292 689 328
rect 694 322 697 338
rect 614 252 617 258
rect 602 238 606 241
rect 606 152 609 158
rect 494 132 497 138
rect 338 88 342 91
rect 494 82 497 88
rect 374 72 377 78
rect 278 63 281 68
rect 242 58 246 61
rect 414 62 417 78
rect 502 62 505 68
rect 510 62 513 148
rect 566 148 574 151
rect 526 142 529 147
rect 574 142 577 148
rect 594 138 598 141
rect 558 132 561 138
rect 614 132 617 228
rect 594 128 598 131
rect 606 128 614 131
rect 526 82 529 128
rect 606 92 609 128
rect 526 72 529 78
rect 474 58 478 61
rect 554 58 558 61
rect 198 52 201 58
rect 368 3 370 7
rect 374 3 377 7
rect 381 3 384 7
rect 566 -18 569 8
rect 566 -22 570 -18
rect 614 -19 618 -18
rect 622 -19 625 258
rect 630 62 633 138
rect 638 92 641 258
rect 646 252 649 288
rect 678 282 681 288
rect 702 272 705 358
rect 710 282 713 368
rect 730 358 734 361
rect 722 348 726 351
rect 670 152 673 168
rect 678 162 681 248
rect 686 192 689 218
rect 682 158 686 161
rect 658 148 662 151
rect 694 92 697 138
rect 658 88 662 91
rect 646 12 649 68
rect 614 -22 625 -19
rect 630 -18 633 8
rect 702 -18 705 268
rect 742 262 745 548
rect 750 462 753 518
rect 750 342 753 368
rect 758 352 761 528
rect 766 472 769 478
rect 782 422 785 548
rect 790 522 793 548
rect 798 492 801 538
rect 806 522 809 748
rect 830 742 833 778
rect 846 752 849 848
rect 814 722 817 738
rect 814 662 817 668
rect 822 592 825 738
rect 830 581 833 738
rect 838 612 841 748
rect 858 718 862 721
rect 846 662 849 708
rect 870 692 873 838
rect 910 752 913 788
rect 918 762 921 858
rect 926 742 929 938
rect 942 881 945 988
rect 958 962 961 1138
rect 966 1132 969 1148
rect 982 1142 985 1258
rect 990 1232 993 1258
rect 1002 1248 1006 1251
rect 1022 1242 1025 1258
rect 994 1168 998 1171
rect 974 1082 977 1118
rect 990 1112 993 1138
rect 982 1072 985 1078
rect 990 1062 993 1098
rect 1014 1072 1017 1118
rect 1038 1092 1041 1248
rect 1126 1162 1129 1168
rect 1142 1152 1145 1238
rect 1286 1232 1289 1258
rect 1294 1232 1297 1258
rect 1334 1242 1337 1268
rect 1342 1262 1345 1268
rect 1374 1262 1377 1348
rect 1390 1282 1393 1318
rect 1406 1272 1409 1318
rect 1422 1292 1425 1528
rect 1458 1518 1462 1521
rect 1502 1492 1505 1668
rect 1518 1482 1521 1618
rect 1470 1472 1473 1478
rect 1526 1472 1529 1518
rect 1542 1472 1545 1528
rect 1550 1482 1553 1518
rect 1558 1502 1561 1588
rect 1566 1522 1569 1668
rect 1594 1658 1598 1661
rect 1666 1658 1670 1661
rect 1730 1658 1734 1661
rect 1646 1612 1649 1618
rect 1654 1612 1657 1658
rect 1686 1642 1689 1658
rect 1702 1652 1705 1658
rect 1590 1560 1593 1579
rect 1574 1552 1577 1558
rect 1558 1482 1561 1498
rect 1574 1492 1577 1548
rect 1582 1492 1585 1538
rect 1622 1532 1625 1538
rect 1638 1522 1641 1528
rect 1678 1522 1681 1618
rect 1710 1562 1713 1658
rect 1726 1562 1729 1618
rect 1614 1482 1617 1508
rect 1638 1482 1641 1518
rect 1718 1512 1721 1518
rect 1734 1502 1737 1548
rect 1570 1468 1574 1471
rect 1446 1452 1449 1458
rect 1442 1348 1446 1351
rect 1470 1342 1473 1468
rect 1486 1452 1489 1458
rect 1494 1432 1497 1468
rect 1646 1462 1649 1488
rect 1702 1482 1705 1488
rect 1686 1462 1689 1468
rect 1546 1458 1550 1461
rect 1566 1452 1569 1458
rect 1486 1362 1489 1378
rect 1430 1282 1433 1328
rect 1478 1292 1481 1308
rect 1486 1272 1489 1318
rect 1510 1312 1513 1338
rect 1518 1292 1521 1328
rect 1506 1288 1510 1291
rect 1498 1278 1502 1281
rect 1470 1262 1473 1268
rect 1534 1262 1537 1338
rect 1542 1332 1545 1418
rect 1598 1382 1601 1458
rect 1630 1392 1633 1448
rect 1654 1422 1657 1450
rect 1742 1422 1745 1658
rect 1750 1592 1753 1668
rect 1770 1658 1774 1661
rect 1790 1582 1793 1618
rect 1798 1592 1801 1658
rect 1566 1352 1569 1368
rect 1638 1362 1641 1378
rect 1574 1342 1577 1348
rect 1598 1342 1601 1358
rect 1630 1352 1633 1358
rect 1610 1348 1617 1351
rect 1598 1322 1601 1328
rect 1550 1262 1553 1318
rect 1358 1252 1361 1258
rect 1214 1152 1217 1158
rect 1326 1152 1329 1158
rect 1334 1152 1337 1228
rect 1050 1148 1054 1151
rect 998 1062 1001 1068
rect 1030 1062 1033 1068
rect 1006 1042 1009 1058
rect 966 992 969 1018
rect 1002 988 1006 991
rect 998 962 1001 968
rect 970 958 974 961
rect 938 878 945 881
rect 958 932 961 938
rect 950 862 953 868
rect 958 862 961 928
rect 966 892 969 938
rect 982 932 985 938
rect 998 902 1001 918
rect 1022 882 1025 1058
rect 1038 891 1041 1018
rect 1046 972 1049 1058
rect 1046 942 1049 948
rect 1054 942 1057 1138
rect 1078 1132 1081 1138
rect 1094 1122 1097 1128
rect 1070 1092 1073 1108
rect 1106 1088 1110 1091
rect 1094 1082 1097 1088
rect 1074 1068 1078 1071
rect 1062 952 1065 1068
rect 1094 1062 1097 1078
rect 1102 952 1105 1018
rect 1126 992 1129 1058
rect 1142 992 1145 1148
rect 1150 1142 1153 1148
rect 1322 1138 1326 1141
rect 1214 1132 1217 1138
rect 1154 1118 1158 1121
rect 1214 1072 1217 1128
rect 1262 1072 1265 1118
rect 1162 1058 1166 1061
rect 1262 1062 1265 1068
rect 1310 1062 1313 1068
rect 1230 1042 1233 1059
rect 1130 948 1134 951
rect 1038 888 1049 891
rect 1014 872 1017 878
rect 990 862 993 868
rect 978 858 982 861
rect 934 842 937 858
rect 950 852 953 858
rect 958 742 961 858
rect 966 792 969 838
rect 974 762 977 778
rect 998 752 1001 858
rect 1006 802 1009 818
rect 1006 792 1009 798
rect 1022 792 1025 858
rect 1030 801 1033 858
rect 1030 798 1041 801
rect 1006 752 1009 768
rect 962 738 966 741
rect 978 738 982 741
rect 888 703 890 707
rect 894 703 897 707
rect 901 703 904 707
rect 926 692 929 738
rect 910 682 913 688
rect 910 672 913 678
rect 858 668 862 671
rect 846 642 849 658
rect 854 652 857 658
rect 862 652 865 658
rect 854 612 857 648
rect 894 622 897 658
rect 838 592 841 598
rect 822 578 833 581
rect 822 542 825 578
rect 918 562 921 648
rect 818 538 822 541
rect 814 462 817 468
rect 814 432 817 448
rect 758 332 761 348
rect 774 342 777 348
rect 758 292 761 318
rect 766 272 769 278
rect 754 268 758 271
rect 774 262 777 328
rect 750 242 753 258
rect 750 152 753 198
rect 782 192 785 418
rect 814 392 817 428
rect 794 378 798 381
rect 806 352 809 388
rect 830 362 833 548
rect 878 538 886 541
rect 878 522 881 538
rect 902 532 905 547
rect 838 462 841 468
rect 878 442 881 518
rect 888 503 890 507
rect 894 503 897 507
rect 901 503 904 507
rect 906 488 910 491
rect 918 462 921 558
rect 950 552 953 708
rect 974 552 977 718
rect 998 712 1001 748
rect 1006 732 1009 738
rect 1026 728 1030 731
rect 1014 692 1017 718
rect 1038 712 1041 798
rect 1046 752 1049 888
rect 1062 882 1065 938
rect 1062 863 1065 868
rect 1142 842 1145 948
rect 1150 942 1153 948
rect 1178 928 1182 931
rect 1150 882 1153 928
rect 1158 892 1161 918
rect 1206 892 1209 1038
rect 1166 862 1169 868
rect 1222 862 1225 948
rect 1262 932 1265 1058
rect 1290 1018 1294 1021
rect 1334 1012 1337 1148
rect 1362 1138 1366 1141
rect 1342 1062 1345 1078
rect 1358 1072 1361 1128
rect 1374 1122 1377 1258
rect 1406 1222 1409 1258
rect 1384 1203 1386 1207
rect 1390 1203 1393 1207
rect 1397 1203 1400 1207
rect 1394 1168 1398 1171
rect 1438 1132 1441 1148
rect 1462 1142 1465 1148
rect 1526 1132 1529 1138
rect 1550 1132 1553 1148
rect 1438 1072 1441 1078
rect 1430 1062 1433 1068
rect 1438 1052 1441 1058
rect 1334 992 1337 1008
rect 1310 960 1313 979
rect 1326 952 1329 958
rect 1238 882 1241 908
rect 1262 901 1265 928
rect 1278 922 1281 938
rect 1262 898 1273 901
rect 1270 882 1273 898
rect 1350 872 1353 1028
rect 1384 1003 1386 1007
rect 1390 1003 1393 1007
rect 1397 1003 1400 1007
rect 1382 962 1385 988
rect 1374 952 1377 958
rect 1358 892 1361 918
rect 1374 862 1377 938
rect 1430 922 1433 938
rect 1446 932 1449 1128
rect 1510 1122 1513 1128
rect 1462 1062 1465 1068
rect 1470 1062 1473 1118
rect 1478 1072 1481 1078
rect 1482 1058 1486 1061
rect 1470 1012 1473 1058
rect 1494 1042 1497 1068
rect 1486 952 1489 958
rect 1406 882 1409 908
rect 1446 882 1449 928
rect 1502 901 1505 1118
rect 1558 1082 1561 1268
rect 1598 1242 1601 1268
rect 1606 1262 1609 1298
rect 1614 1272 1617 1348
rect 1630 1272 1633 1278
rect 1638 1272 1641 1358
rect 1662 1352 1665 1358
rect 1686 1352 1689 1368
rect 1674 1348 1678 1351
rect 1670 1332 1673 1338
rect 1646 1262 1649 1278
rect 1670 1262 1673 1278
rect 1650 1258 1654 1261
rect 1622 1252 1625 1258
rect 1598 1162 1601 1238
rect 1610 1178 1614 1181
rect 1622 1152 1625 1208
rect 1610 1148 1614 1151
rect 1526 912 1529 918
rect 1502 898 1510 901
rect 1478 872 1481 888
rect 1494 872 1497 878
rect 1534 862 1537 958
rect 1550 952 1553 1058
rect 1558 992 1561 1059
rect 1574 952 1577 1098
rect 1614 1092 1617 1138
rect 1622 1102 1625 1148
rect 1630 1142 1633 1258
rect 1662 1252 1665 1258
rect 1670 1212 1673 1258
rect 1634 1128 1638 1131
rect 1646 1092 1649 1128
rect 1622 1081 1625 1088
rect 1614 1078 1625 1081
rect 1590 1002 1593 1068
rect 1598 1052 1601 1058
rect 1614 1052 1617 1078
rect 1654 1072 1657 1158
rect 1670 1142 1673 1178
rect 1678 1092 1681 1328
rect 1686 1262 1689 1268
rect 1686 1131 1689 1218
rect 1694 1182 1697 1318
rect 1702 1282 1705 1418
rect 1742 1392 1745 1408
rect 1734 1352 1737 1388
rect 1710 1322 1713 1348
rect 1726 1342 1729 1348
rect 1734 1282 1737 1348
rect 1750 1272 1753 1478
rect 1758 1372 1761 1518
rect 1758 1352 1761 1358
rect 1766 1282 1769 1528
rect 1774 1512 1777 1548
rect 1778 1418 1782 1421
rect 1782 1352 1785 1358
rect 1782 1332 1785 1338
rect 1694 1152 1697 1158
rect 1710 1152 1713 1168
rect 1718 1161 1721 1258
rect 1734 1252 1737 1259
rect 1718 1158 1726 1161
rect 1686 1128 1697 1131
rect 1686 1092 1689 1118
rect 1694 1081 1697 1128
rect 1690 1078 1697 1081
rect 1702 1072 1705 1138
rect 1626 1068 1630 1071
rect 1666 1068 1670 1071
rect 1626 1058 1630 1061
rect 1630 1022 1633 1058
rect 1598 952 1601 988
rect 1606 962 1609 968
rect 1630 952 1633 1008
rect 1638 952 1641 1068
rect 1646 1062 1649 1068
rect 1654 1052 1657 1068
rect 1642 948 1646 951
rect 1582 942 1585 948
rect 1622 942 1625 948
rect 1630 892 1633 948
rect 1610 888 1614 891
rect 1578 878 1582 881
rect 1638 872 1641 878
rect 1646 872 1649 918
rect 1594 868 1598 871
rect 1654 862 1657 1018
rect 1662 922 1665 1058
rect 1670 911 1673 1048
rect 1670 908 1681 911
rect 1670 882 1673 888
rect 1678 872 1681 908
rect 1686 872 1689 1068
rect 1698 1058 1702 1061
rect 1710 952 1713 958
rect 1206 858 1214 861
rect 1226 858 1230 861
rect 1594 858 1601 861
rect 1174 852 1177 858
rect 1190 852 1193 858
rect 1142 792 1145 818
rect 1158 792 1161 848
rect 1206 812 1209 858
rect 1234 848 1238 851
rect 1054 752 1057 778
rect 1086 752 1089 778
rect 1110 752 1113 788
rect 1138 778 1142 781
rect 1126 768 1134 771
rect 1126 762 1129 768
rect 1182 752 1185 768
rect 1066 748 1070 751
rect 982 682 985 688
rect 982 663 985 668
rect 946 548 950 551
rect 962 538 966 541
rect 982 532 985 598
rect 998 552 1001 688
rect 1014 672 1017 678
rect 1034 668 1038 671
rect 1006 592 1009 598
rect 970 528 974 531
rect 974 482 977 488
rect 978 478 982 481
rect 990 481 993 548
rect 998 542 1001 548
rect 1006 492 1009 578
rect 990 478 1001 481
rect 926 462 929 478
rect 934 472 937 478
rect 978 458 982 461
rect 838 362 841 368
rect 826 348 830 351
rect 798 332 801 348
rect 818 328 822 331
rect 790 162 793 318
rect 798 292 801 328
rect 826 288 830 291
rect 810 278 814 281
rect 798 262 801 268
rect 802 188 806 191
rect 718 142 721 148
rect 738 138 742 141
rect 814 141 817 278
rect 806 138 817 141
rect 718 63 721 68
rect 734 62 737 118
rect 782 72 785 78
rect 778 58 782 61
rect 790 12 793 138
rect 774 -18 777 8
rect 806 -18 809 138
rect 830 72 833 138
rect 838 92 841 338
rect 854 322 857 338
rect 870 332 873 348
rect 878 342 881 438
rect 886 352 889 368
rect 894 352 897 438
rect 918 372 921 458
rect 910 352 913 358
rect 878 272 881 338
rect 888 303 890 307
rect 894 303 897 307
rect 901 303 904 307
rect 926 292 929 458
rect 990 392 993 468
rect 942 332 945 388
rect 974 351 977 358
rect 958 342 961 348
rect 918 282 921 288
rect 954 268 958 271
rect 878 172 881 268
rect 886 263 889 268
rect 998 262 1001 478
rect 1014 472 1017 478
rect 1006 432 1009 468
rect 1030 462 1033 508
rect 1038 492 1041 628
rect 1046 482 1049 728
rect 1054 652 1057 748
rect 1130 738 1142 741
rect 1162 738 1182 741
rect 1062 662 1065 738
rect 1102 722 1105 738
rect 1078 692 1081 718
rect 1102 682 1105 698
rect 1158 691 1161 728
rect 1190 722 1193 728
rect 1182 692 1185 708
rect 1158 688 1166 691
rect 1070 662 1073 668
rect 1110 662 1113 688
rect 1170 678 1174 681
rect 1062 642 1065 658
rect 1066 547 1070 550
rect 1054 522 1057 538
rect 1102 532 1105 598
rect 1150 552 1153 568
rect 1158 552 1161 648
rect 1174 592 1177 668
rect 1206 662 1209 808
rect 1238 782 1241 848
rect 1222 752 1225 778
rect 1234 768 1238 771
rect 1214 682 1217 738
rect 1238 712 1241 748
rect 1246 742 1249 768
rect 1254 752 1257 858
rect 1278 812 1281 858
rect 1330 818 1334 821
rect 1286 752 1289 768
rect 1266 748 1270 751
rect 1214 672 1217 678
rect 1230 662 1233 668
rect 1238 662 1241 668
rect 1186 658 1190 661
rect 1198 652 1201 658
rect 1146 548 1150 551
rect 1118 542 1121 548
rect 1182 542 1185 588
rect 1190 582 1193 588
rect 1206 552 1209 658
rect 1214 592 1217 618
rect 1238 552 1241 598
rect 1078 482 1081 498
rect 1090 488 1094 491
rect 1026 458 1030 461
rect 1014 402 1017 458
rect 1046 432 1049 468
rect 1034 388 1038 391
rect 1006 292 1009 358
rect 1046 332 1049 368
rect 1042 328 1046 331
rect 1006 262 1009 288
rect 1054 282 1057 458
rect 1062 382 1065 468
rect 1070 352 1073 418
rect 1062 342 1065 348
rect 1086 342 1089 478
rect 1102 472 1105 518
rect 1166 512 1169 528
rect 1182 492 1185 498
rect 1190 492 1193 548
rect 1242 538 1246 541
rect 1126 462 1129 468
rect 1206 462 1209 478
rect 1214 472 1217 488
rect 1222 482 1225 498
rect 1238 472 1241 488
rect 1242 458 1246 461
rect 1186 448 1190 451
rect 1098 368 1102 371
rect 1078 322 1081 328
rect 1038 262 1041 268
rect 978 258 982 261
rect 998 212 1001 258
rect 862 151 865 158
rect 878 142 881 168
rect 910 132 913 188
rect 958 152 961 158
rect 966 152 969 208
rect 978 188 982 191
rect 1006 152 1009 168
rect 1038 151 1041 158
rect 926 142 929 148
rect 888 103 890 107
rect 894 103 897 107
rect 901 103 904 107
rect 950 92 953 148
rect 1070 132 1073 188
rect 1078 121 1081 308
rect 1094 152 1097 348
rect 1142 332 1145 348
rect 1142 262 1145 268
rect 1158 262 1161 338
rect 1166 292 1169 448
rect 1206 392 1209 448
rect 1222 362 1225 458
rect 1254 392 1257 748
rect 1294 742 1297 748
rect 1310 732 1313 768
rect 1270 682 1273 698
rect 1270 652 1273 659
rect 1262 492 1265 528
rect 1274 518 1278 521
rect 1274 468 1278 471
rect 1302 462 1305 548
rect 1310 472 1313 608
rect 1318 482 1321 818
rect 1334 792 1337 808
rect 1326 752 1329 758
rect 1326 732 1329 748
rect 1342 722 1345 858
rect 1374 852 1377 858
rect 1446 822 1449 850
rect 1384 803 1386 807
rect 1390 803 1393 807
rect 1397 803 1400 807
rect 1350 752 1353 758
rect 1358 752 1361 798
rect 1534 791 1537 858
rect 1534 788 1545 791
rect 1378 768 1382 771
rect 1358 672 1361 678
rect 1342 662 1345 668
rect 1346 658 1350 661
rect 1362 658 1366 661
rect 1374 632 1377 748
rect 1382 662 1385 708
rect 1390 672 1393 778
rect 1510 760 1513 779
rect 1542 752 1545 788
rect 1434 748 1438 751
rect 1414 672 1417 688
rect 1422 662 1425 748
rect 1446 711 1449 728
rect 1446 708 1457 711
rect 1438 662 1441 678
rect 1382 621 1385 658
rect 1374 618 1385 621
rect 1366 602 1369 618
rect 1326 492 1329 578
rect 1334 551 1337 558
rect 1350 542 1353 548
rect 1366 522 1369 528
rect 1310 462 1313 468
rect 1334 462 1337 468
rect 1342 462 1345 468
rect 1366 462 1369 478
rect 1274 458 1278 461
rect 1222 352 1225 358
rect 1202 348 1206 351
rect 1202 338 1206 341
rect 1226 328 1230 331
rect 1238 312 1241 338
rect 1254 312 1257 318
rect 1262 301 1265 448
rect 1254 298 1265 301
rect 1270 322 1273 338
rect 1254 292 1257 298
rect 1114 258 1118 261
rect 1162 248 1166 251
rect 1102 162 1105 168
rect 1118 152 1121 198
rect 1126 152 1129 208
rect 1174 162 1177 268
rect 1190 262 1193 288
rect 1242 278 1246 281
rect 1262 272 1265 278
rect 1218 268 1222 271
rect 1270 262 1273 318
rect 1302 292 1305 458
rect 1326 412 1329 448
rect 1326 342 1329 408
rect 1358 351 1361 418
rect 1342 332 1345 338
rect 1366 292 1369 438
rect 1374 322 1377 618
rect 1384 603 1386 607
rect 1390 603 1393 607
rect 1397 603 1400 607
rect 1422 582 1425 658
rect 1434 648 1438 651
rect 1446 622 1449 668
rect 1430 562 1433 618
rect 1386 558 1390 561
rect 1430 552 1433 558
rect 1438 552 1441 558
rect 1410 548 1414 551
rect 1382 542 1385 548
rect 1422 492 1425 538
rect 1438 512 1441 548
rect 1454 542 1457 708
rect 1470 692 1473 718
rect 1542 711 1545 738
rect 1558 722 1561 728
rect 1534 708 1545 711
rect 1534 692 1537 708
rect 1542 682 1545 688
rect 1518 678 1537 681
rect 1462 642 1465 678
rect 1518 672 1521 678
rect 1482 668 1502 671
rect 1534 671 1537 678
rect 1534 668 1542 671
rect 1478 652 1481 658
rect 1518 602 1521 658
rect 1526 652 1529 668
rect 1550 652 1553 698
rect 1478 552 1481 578
rect 1454 532 1457 538
rect 1384 403 1386 407
rect 1390 403 1393 407
rect 1397 403 1400 407
rect 1406 392 1409 478
rect 1462 392 1465 478
rect 1478 452 1481 468
rect 1494 462 1497 568
rect 1542 552 1545 628
rect 1574 592 1577 668
rect 1574 552 1577 568
rect 1554 548 1558 551
rect 1502 462 1505 538
rect 1542 522 1545 548
rect 1534 512 1537 518
rect 1486 422 1489 458
rect 1418 388 1422 391
rect 1494 391 1497 458
rect 1486 388 1497 391
rect 1422 358 1430 361
rect 1390 272 1393 318
rect 1422 292 1425 358
rect 1326 262 1329 268
rect 1182 212 1185 258
rect 1138 158 1142 161
rect 1158 152 1161 158
rect 1178 148 1182 151
rect 1190 151 1193 258
rect 1242 248 1246 251
rect 1214 152 1217 208
rect 1222 152 1225 158
rect 1186 148 1193 151
rect 1202 148 1206 151
rect 1242 148 1246 151
rect 1150 142 1153 148
rect 1270 142 1273 258
rect 1302 252 1305 258
rect 1366 242 1369 248
rect 1366 192 1369 218
rect 1298 148 1302 151
rect 1194 128 1198 131
rect 1070 118 1081 121
rect 966 92 969 98
rect 1070 92 1073 118
rect 1046 72 1049 88
rect 1118 72 1121 88
rect 862 62 865 68
rect 902 62 905 68
rect 930 58 934 61
rect 894 52 897 58
rect 958 12 961 68
rect 1026 59 1030 62
rect 1078 42 1081 68
rect 1126 62 1129 118
rect 1134 102 1137 128
rect 1166 62 1169 118
rect 1174 92 1177 128
rect 1234 118 1238 121
rect 1230 92 1233 108
rect 1270 92 1273 138
rect 1366 92 1369 168
rect 1226 78 1230 81
rect 942 -18 945 8
rect 630 -22 634 -18
rect 702 -22 706 -18
rect 774 -22 778 -18
rect 806 -22 810 -18
rect 942 -22 946 -18
rect 1062 -19 1065 38
rect 1070 -19 1074 -18
rect 1062 -22 1074 -19
rect 1078 -19 1081 38
rect 1198 -18 1201 78
rect 1214 72 1217 78
rect 1218 58 1222 61
rect 1086 -19 1090 -18
rect 1078 -22 1090 -19
rect 1198 -22 1202 -18
rect 1246 -19 1250 -18
rect 1254 -19 1257 78
rect 1270 72 1273 88
rect 1294 62 1297 78
rect 1358 72 1361 78
rect 1374 52 1377 228
rect 1384 203 1386 207
rect 1390 203 1393 207
rect 1397 203 1400 207
rect 1406 182 1409 258
rect 1414 232 1417 248
rect 1406 152 1409 168
rect 1430 152 1433 308
rect 1450 288 1454 291
rect 1438 282 1441 288
rect 1462 281 1465 348
rect 1470 322 1473 338
rect 1454 278 1465 281
rect 1454 222 1457 278
rect 1446 152 1449 218
rect 1462 192 1465 248
rect 1486 172 1489 388
rect 1502 342 1505 458
rect 1510 352 1513 418
rect 1518 402 1521 458
rect 1534 322 1537 468
rect 1542 452 1545 458
rect 1534 272 1537 318
rect 1550 282 1553 508
rect 1558 492 1561 538
rect 1566 512 1569 518
rect 1566 492 1569 498
rect 1562 448 1569 451
rect 1558 292 1561 438
rect 1566 292 1569 448
rect 1582 442 1585 658
rect 1598 642 1601 858
rect 1646 858 1654 861
rect 1622 852 1625 858
rect 1622 662 1625 748
rect 1638 712 1641 718
rect 1630 672 1633 678
rect 1638 662 1641 688
rect 1646 662 1649 858
rect 1670 842 1673 858
rect 1654 752 1657 758
rect 1662 742 1665 748
rect 1670 682 1673 688
rect 1678 672 1681 868
rect 1686 862 1689 868
rect 1710 862 1713 878
rect 1698 858 1702 861
rect 1694 752 1697 858
rect 1718 852 1721 1158
rect 1734 1132 1737 1148
rect 1742 1112 1745 1128
rect 1750 1122 1753 1218
rect 1766 1072 1769 1258
rect 1762 1058 1766 1061
rect 1726 991 1729 1038
rect 1766 992 1769 1048
rect 1790 992 1793 1568
rect 1798 1242 1801 1328
rect 1798 1212 1801 1218
rect 1726 988 1737 991
rect 1734 942 1737 988
rect 1750 932 1753 948
rect 1734 892 1737 918
rect 1774 912 1777 948
rect 1798 892 1801 1038
rect 1730 878 1734 881
rect 1782 862 1785 868
rect 1706 848 1710 851
rect 1706 788 1710 791
rect 1754 748 1758 751
rect 1686 742 1689 748
rect 1686 682 1689 718
rect 1758 682 1761 738
rect 1798 692 1801 878
rect 1610 658 1614 661
rect 1650 658 1654 661
rect 1598 582 1601 618
rect 1614 552 1617 598
rect 1610 538 1614 541
rect 1598 482 1601 528
rect 1598 462 1601 468
rect 1614 462 1617 508
rect 1622 422 1625 658
rect 1630 561 1633 638
rect 1638 602 1641 618
rect 1654 552 1657 558
rect 1662 552 1665 668
rect 1730 658 1734 661
rect 1670 652 1673 658
rect 1678 592 1681 658
rect 1698 618 1702 621
rect 1686 552 1689 568
rect 1662 492 1665 548
rect 1686 492 1689 538
rect 1694 492 1697 608
rect 1706 588 1710 591
rect 1702 482 1705 558
rect 1742 552 1745 668
rect 1790 582 1793 678
rect 1662 472 1665 478
rect 1582 392 1585 398
rect 1618 348 1622 351
rect 1582 328 1590 331
rect 1582 272 1585 328
rect 1590 322 1593 328
rect 1498 258 1502 261
rect 1510 252 1513 258
rect 1566 232 1569 248
rect 1470 152 1473 168
rect 1486 152 1489 158
rect 1526 152 1529 178
rect 1558 151 1561 158
rect 1582 152 1585 258
rect 1590 182 1593 218
rect 1598 192 1601 278
rect 1614 262 1617 268
rect 1382 142 1385 148
rect 1478 142 1481 148
rect 1382 82 1385 88
rect 1398 78 1406 81
rect 1398 72 1401 78
rect 1446 62 1449 128
rect 1462 72 1465 138
rect 1494 132 1497 148
rect 1518 142 1521 148
rect 1542 72 1545 138
rect 1602 88 1606 91
rect 1614 72 1617 258
rect 1622 192 1625 198
rect 1630 152 1633 408
rect 1638 352 1641 358
rect 1646 352 1649 408
rect 1670 402 1673 458
rect 1686 452 1689 468
rect 1742 462 1745 548
rect 1766 542 1769 547
rect 1694 452 1697 458
rect 1742 452 1745 458
rect 1694 352 1697 448
rect 1714 418 1718 421
rect 1706 348 1710 351
rect 1650 318 1654 321
rect 1694 302 1697 348
rect 1702 292 1705 338
rect 1694 282 1697 288
rect 1710 282 1713 328
rect 1718 292 1721 398
rect 1750 352 1753 518
rect 1762 458 1766 461
rect 1766 392 1769 438
rect 1758 352 1761 358
rect 1774 292 1777 508
rect 1798 491 1801 618
rect 1790 488 1801 491
rect 1782 352 1785 368
rect 1738 268 1742 271
rect 1790 262 1793 488
rect 1798 272 1801 288
rect 1738 258 1742 261
rect 1646 192 1649 258
rect 1718 242 1721 248
rect 1686 192 1689 238
rect 1694 222 1697 228
rect 1694 162 1697 218
rect 1734 192 1737 248
rect 1706 158 1710 161
rect 1722 158 1726 161
rect 1662 152 1665 158
rect 1642 148 1646 151
rect 1630 142 1633 148
rect 1498 68 1502 71
rect 1462 62 1465 68
rect 1534 63 1537 68
rect 1442 58 1446 61
rect 1498 58 1502 61
rect 1638 62 1641 108
rect 1678 92 1681 138
rect 1742 132 1745 228
rect 1758 162 1761 258
rect 1782 222 1785 248
rect 1758 152 1761 158
rect 1790 152 1793 168
rect 1778 148 1782 151
rect 1706 128 1710 131
rect 1718 102 1721 128
rect 1766 112 1769 118
rect 1694 92 1697 98
rect 1790 92 1793 98
rect 1710 72 1713 78
rect 1726 63 1729 68
rect 1470 52 1473 58
rect 1384 3 1386 7
rect 1390 3 1393 7
rect 1397 3 1400 7
rect 1246 -22 1257 -19
<< m3contact >>
rect 14 1688 18 1692
rect 150 1688 154 1692
rect 318 1688 322 1692
rect 430 1688 434 1692
rect 518 1688 522 1692
rect 62 1668 66 1672
rect 38 1658 42 1662
rect 94 1648 98 1652
rect 150 1618 154 1622
rect 62 1608 66 1612
rect 126 1608 130 1612
rect 54 1548 58 1552
rect 38 1538 42 1542
rect 222 1608 226 1612
rect 190 1558 194 1562
rect 206 1548 210 1552
rect 222 1548 226 1552
rect 126 1538 130 1542
rect 110 1528 114 1532
rect 94 1478 98 1482
rect 110 1478 114 1482
rect 118 1468 122 1472
rect 134 1468 138 1472
rect 158 1538 162 1542
rect 190 1538 194 1542
rect 166 1528 170 1532
rect 158 1478 162 1482
rect 46 1458 50 1462
rect 126 1458 130 1462
rect 198 1478 202 1482
rect 286 1608 290 1612
rect 262 1588 266 1592
rect 262 1558 266 1562
rect 254 1458 258 1462
rect 190 1448 194 1452
rect 174 1438 178 1442
rect 198 1368 202 1372
rect 150 1358 154 1362
rect 206 1358 210 1362
rect 110 1348 114 1352
rect 142 1348 146 1352
rect 62 1338 66 1342
rect 46 1318 50 1322
rect 62 1308 66 1312
rect 94 1308 98 1312
rect 198 1318 202 1322
rect 118 1278 122 1282
rect 22 1258 26 1262
rect 54 1258 58 1262
rect 110 1258 114 1262
rect 38 1248 42 1252
rect 46 1238 50 1242
rect 22 1168 26 1172
rect 38 1158 42 1162
rect 70 1188 74 1192
rect 102 1248 106 1252
rect 94 1168 98 1172
rect 78 1158 82 1162
rect 22 1148 26 1152
rect 54 1148 58 1152
rect 38 1048 42 1052
rect 30 948 34 952
rect 30 858 34 862
rect 30 748 34 752
rect 38 728 42 732
rect 6 648 10 652
rect 22 548 26 552
rect 62 1138 66 1142
rect 62 1088 66 1092
rect 286 1448 290 1452
rect 270 1378 274 1382
rect 254 1368 258 1372
rect 262 1368 266 1372
rect 222 1358 226 1362
rect 230 1348 234 1352
rect 238 1348 242 1352
rect 230 1308 234 1312
rect 222 1278 226 1282
rect 342 1678 346 1682
rect 890 1703 894 1707
rect 897 1703 901 1707
rect 1254 1688 1258 1692
rect 702 1678 706 1682
rect 718 1678 722 1682
rect 814 1678 818 1682
rect 830 1678 834 1682
rect 854 1678 858 1682
rect 870 1678 874 1682
rect 422 1668 426 1672
rect 494 1668 498 1672
rect 366 1658 370 1662
rect 414 1658 418 1662
rect 382 1638 386 1642
rect 342 1628 346 1632
rect 326 1578 330 1582
rect 370 1603 374 1607
rect 377 1603 381 1607
rect 542 1658 546 1662
rect 462 1648 466 1652
rect 614 1658 618 1662
rect 598 1628 602 1632
rect 574 1588 578 1592
rect 638 1588 642 1592
rect 542 1578 546 1582
rect 398 1518 402 1522
rect 478 1538 482 1542
rect 494 1538 498 1542
rect 422 1498 426 1502
rect 430 1498 434 1502
rect 406 1468 410 1472
rect 422 1468 426 1472
rect 326 1458 330 1462
rect 390 1458 394 1462
rect 422 1448 426 1452
rect 390 1428 394 1432
rect 422 1428 426 1432
rect 370 1403 374 1407
rect 377 1403 381 1407
rect 406 1388 410 1392
rect 366 1378 370 1382
rect 342 1368 346 1372
rect 278 1358 282 1362
rect 294 1358 298 1362
rect 302 1358 306 1362
rect 278 1348 282 1352
rect 334 1348 338 1352
rect 310 1338 314 1342
rect 358 1338 362 1342
rect 390 1328 394 1332
rect 374 1318 378 1322
rect 158 1248 162 1252
rect 214 1248 218 1252
rect 166 1158 170 1162
rect 158 1148 162 1152
rect 182 1138 186 1142
rect 198 1138 202 1142
rect 158 1128 162 1132
rect 126 1088 130 1092
rect 166 1088 170 1092
rect 118 1068 122 1072
rect 134 1068 138 1072
rect 126 1058 130 1062
rect 94 1028 98 1032
rect 94 978 98 982
rect 358 1288 362 1292
rect 350 1278 354 1282
rect 294 1268 298 1272
rect 254 1238 258 1242
rect 254 1178 258 1182
rect 318 1158 322 1162
rect 390 1268 394 1272
rect 390 1258 394 1262
rect 398 1228 402 1232
rect 374 1218 378 1222
rect 370 1203 374 1207
rect 377 1203 381 1207
rect 398 1178 402 1182
rect 366 1148 370 1152
rect 326 1138 330 1142
rect 350 1138 354 1142
rect 254 1128 258 1132
rect 230 1118 234 1122
rect 206 1078 210 1082
rect 198 1068 202 1072
rect 150 1018 154 1022
rect 134 978 138 982
rect 158 988 162 992
rect 150 958 154 962
rect 182 978 186 982
rect 198 978 202 982
rect 166 958 170 962
rect 118 948 122 952
rect 126 948 130 952
rect 142 948 146 952
rect 102 938 106 942
rect 118 898 122 902
rect 102 888 106 892
rect 110 878 114 882
rect 150 888 154 892
rect 214 948 218 952
rect 206 928 210 932
rect 142 878 146 882
rect 174 878 178 882
rect 102 858 106 862
rect 174 858 178 862
rect 182 848 186 852
rect 94 738 98 742
rect 126 778 130 782
rect 118 728 122 732
rect 62 718 66 722
rect 86 698 90 702
rect 102 698 106 702
rect 54 668 58 672
rect 102 688 106 692
rect 110 688 114 692
rect 78 658 82 662
rect 94 588 98 592
rect 46 568 50 572
rect 70 558 74 562
rect 54 548 58 552
rect 30 538 34 542
rect 158 748 162 752
rect 142 738 146 742
rect 150 728 154 732
rect 158 718 162 722
rect 222 918 226 922
rect 214 898 218 902
rect 206 878 210 882
rect 198 868 202 872
rect 222 868 226 872
rect 310 1108 314 1112
rect 342 1128 346 1132
rect 366 1118 370 1122
rect 246 1088 250 1092
rect 302 1088 306 1092
rect 278 1078 282 1082
rect 238 958 242 962
rect 246 948 250 952
rect 254 938 258 942
rect 246 928 250 932
rect 254 918 258 922
rect 254 888 258 892
rect 278 1038 282 1042
rect 270 878 274 882
rect 262 858 266 862
rect 302 958 306 962
rect 294 948 298 952
rect 286 888 290 892
rect 294 868 298 872
rect 278 848 282 852
rect 214 838 218 842
rect 198 778 202 782
rect 222 778 226 782
rect 190 758 194 762
rect 238 838 242 842
rect 254 838 258 842
rect 302 838 306 842
rect 278 828 282 832
rect 262 788 266 792
rect 238 768 242 772
rect 214 758 218 762
rect 230 748 234 752
rect 302 748 306 752
rect 390 1088 394 1092
rect 414 1218 418 1222
rect 326 1048 330 1052
rect 326 1018 330 1022
rect 318 928 322 932
rect 370 1003 374 1007
rect 377 1003 381 1007
rect 358 968 362 972
rect 382 968 386 972
rect 366 958 370 962
rect 334 858 338 862
rect 350 858 354 862
rect 374 908 378 912
rect 350 838 354 842
rect 390 838 394 842
rect 438 1488 442 1492
rect 502 1518 506 1522
rect 518 1528 522 1532
rect 510 1508 514 1512
rect 494 1498 498 1502
rect 518 1498 522 1502
rect 478 1468 482 1472
rect 494 1468 498 1472
rect 462 1438 466 1442
rect 430 1328 434 1332
rect 430 1288 434 1292
rect 606 1558 610 1562
rect 878 1658 882 1662
rect 806 1648 810 1652
rect 1022 1658 1026 1662
rect 1046 1658 1050 1662
rect 1110 1658 1114 1662
rect 918 1648 922 1652
rect 942 1648 946 1652
rect 878 1638 882 1642
rect 1006 1638 1010 1642
rect 742 1628 746 1632
rect 726 1618 730 1622
rect 694 1608 698 1612
rect 726 1578 730 1582
rect 702 1558 706 1562
rect 806 1558 810 1562
rect 598 1548 602 1552
rect 678 1548 682 1552
rect 790 1548 794 1552
rect 566 1488 570 1492
rect 526 1458 530 1462
rect 542 1458 546 1462
rect 830 1547 834 1551
rect 638 1538 642 1542
rect 726 1538 730 1542
rect 766 1538 770 1542
rect 734 1528 738 1532
rect 614 1508 618 1512
rect 598 1488 602 1492
rect 622 1478 626 1482
rect 646 1478 650 1482
rect 630 1468 634 1472
rect 662 1468 666 1472
rect 606 1448 610 1452
rect 654 1448 658 1452
rect 606 1418 610 1422
rect 558 1368 562 1372
rect 654 1378 658 1382
rect 614 1368 618 1372
rect 662 1368 666 1372
rect 582 1358 586 1362
rect 590 1358 594 1362
rect 478 1348 482 1352
rect 502 1348 506 1352
rect 534 1348 538 1352
rect 518 1338 522 1342
rect 526 1328 530 1332
rect 494 1318 498 1322
rect 446 1308 450 1312
rect 454 1308 458 1312
rect 438 1268 442 1272
rect 510 1298 514 1302
rect 534 1278 538 1282
rect 454 1268 458 1272
rect 534 1268 538 1272
rect 438 1248 442 1252
rect 430 1168 434 1172
rect 502 1168 506 1172
rect 446 1158 450 1162
rect 470 1148 474 1152
rect 422 1138 426 1142
rect 542 1258 546 1262
rect 518 1218 522 1222
rect 422 1128 426 1132
rect 558 1338 562 1342
rect 734 1508 738 1512
rect 686 1428 690 1432
rect 686 1408 690 1412
rect 702 1388 706 1392
rect 718 1358 722 1362
rect 806 1498 810 1502
rect 774 1388 778 1392
rect 758 1358 762 1362
rect 934 1588 938 1592
rect 902 1548 906 1552
rect 918 1548 922 1552
rect 1254 1648 1258 1652
rect 1174 1588 1178 1592
rect 1054 1568 1058 1572
rect 1070 1568 1074 1572
rect 1126 1568 1130 1572
rect 1142 1568 1146 1572
rect 1014 1558 1018 1562
rect 1014 1548 1018 1552
rect 918 1528 922 1532
rect 1006 1528 1010 1532
rect 966 1518 970 1522
rect 974 1518 978 1522
rect 822 1458 826 1462
rect 838 1458 842 1462
rect 846 1458 850 1462
rect 890 1503 894 1507
rect 897 1503 901 1507
rect 982 1498 986 1502
rect 926 1468 930 1472
rect 934 1458 938 1462
rect 990 1488 994 1492
rect 1030 1538 1034 1542
rect 1038 1518 1042 1522
rect 1046 1518 1050 1522
rect 1014 1498 1018 1502
rect 1022 1498 1026 1502
rect 1014 1478 1018 1482
rect 998 1458 1002 1462
rect 798 1448 802 1452
rect 814 1448 818 1452
rect 878 1448 882 1452
rect 806 1428 810 1432
rect 790 1418 794 1422
rect 782 1348 786 1352
rect 726 1338 730 1342
rect 614 1328 618 1332
rect 582 1318 586 1322
rect 590 1298 594 1302
rect 606 1268 610 1272
rect 614 1268 618 1272
rect 598 1258 602 1262
rect 606 1258 610 1262
rect 678 1328 682 1332
rect 710 1328 714 1332
rect 798 1378 802 1382
rect 734 1318 738 1322
rect 638 1298 642 1302
rect 630 1288 634 1292
rect 638 1268 642 1272
rect 670 1298 674 1302
rect 702 1298 706 1302
rect 678 1268 682 1272
rect 686 1268 690 1272
rect 662 1258 666 1262
rect 646 1248 650 1252
rect 758 1288 762 1292
rect 726 1258 730 1262
rect 718 1248 722 1252
rect 742 1248 746 1252
rect 638 1238 642 1242
rect 662 1238 666 1242
rect 606 1228 610 1232
rect 726 1228 730 1232
rect 718 1168 722 1172
rect 878 1418 882 1422
rect 934 1418 938 1422
rect 926 1358 930 1362
rect 854 1348 858 1352
rect 870 1348 874 1352
rect 926 1348 930 1352
rect 822 1328 826 1332
rect 790 1258 794 1262
rect 774 1248 778 1252
rect 766 1218 770 1222
rect 742 1168 746 1172
rect 566 1148 570 1152
rect 710 1148 714 1152
rect 470 1118 474 1122
rect 462 1088 466 1092
rect 542 1098 546 1102
rect 654 1128 658 1132
rect 694 1128 698 1132
rect 598 1108 602 1112
rect 630 1108 634 1112
rect 550 1078 554 1082
rect 558 1078 562 1082
rect 574 1078 578 1082
rect 414 1068 418 1072
rect 462 1068 466 1072
rect 526 1068 530 1072
rect 574 1068 578 1072
rect 422 1058 426 1062
rect 478 1048 482 1052
rect 406 1038 410 1042
rect 430 1038 434 1042
rect 510 1048 514 1052
rect 510 1038 514 1042
rect 486 1028 490 1032
rect 494 1028 498 1032
rect 510 1028 514 1032
rect 478 1008 482 1012
rect 454 998 458 1002
rect 406 978 410 982
rect 462 978 466 982
rect 502 978 506 982
rect 422 948 426 952
rect 486 968 490 972
rect 478 958 482 962
rect 470 948 474 952
rect 422 938 426 942
rect 446 938 450 942
rect 462 938 466 942
rect 406 918 410 922
rect 430 928 434 932
rect 454 928 458 932
rect 478 888 482 892
rect 438 868 442 872
rect 446 858 450 862
rect 406 848 410 852
rect 398 818 402 822
rect 370 803 374 807
rect 377 803 381 807
rect 390 798 394 802
rect 390 778 394 782
rect 374 748 378 752
rect 182 688 186 692
rect 206 728 210 732
rect 286 688 290 692
rect 254 678 258 682
rect 262 678 266 682
rect 278 678 282 682
rect 286 678 290 682
rect 198 668 202 672
rect 222 668 226 672
rect 262 668 266 672
rect 142 658 146 662
rect 134 558 138 562
rect 214 658 218 662
rect 238 658 242 662
rect 190 648 194 652
rect 198 648 202 652
rect 190 638 194 642
rect 62 528 66 532
rect 78 488 82 492
rect 94 498 98 502
rect 166 528 170 532
rect 174 508 178 512
rect 206 588 210 592
rect 238 588 242 592
rect 222 568 226 572
rect 278 568 282 572
rect 246 558 250 562
rect 222 548 226 552
rect 326 658 330 662
rect 382 658 386 662
rect 262 548 266 552
rect 286 548 290 552
rect 302 548 306 552
rect 246 538 250 542
rect 214 528 218 532
rect 198 508 202 512
rect 166 478 170 482
rect 86 448 90 452
rect 126 468 130 472
rect 166 458 170 462
rect 150 438 154 442
rect 38 358 42 362
rect 142 398 146 402
rect 134 358 138 362
rect 190 448 194 452
rect 230 458 234 462
rect 206 428 210 432
rect 206 398 210 402
rect 182 358 186 362
rect 46 348 50 352
rect 102 348 106 352
rect 94 298 98 302
rect 62 288 66 292
rect 126 268 130 272
rect 46 258 50 262
rect 118 258 122 262
rect 38 248 42 252
rect 14 158 18 162
rect 222 338 226 342
rect 190 318 194 322
rect 174 298 178 302
rect 182 288 186 292
rect 214 288 218 292
rect 158 278 162 282
rect 174 278 178 282
rect 150 268 154 272
rect 158 268 162 272
rect 134 248 138 252
rect 150 248 154 252
rect 94 178 98 182
rect 46 168 50 172
rect 54 158 58 162
rect 38 148 42 152
rect 62 148 66 152
rect 78 148 82 152
rect 62 88 66 92
rect 54 68 58 72
rect 110 148 114 152
rect 126 128 130 132
rect 94 98 98 102
rect 110 78 114 82
rect 254 438 258 442
rect 206 258 210 262
rect 190 178 194 182
rect 230 248 234 252
rect 222 168 226 172
rect 206 148 210 152
rect 222 148 226 152
rect 166 128 170 132
rect 190 118 194 122
rect 198 108 202 112
rect 166 98 170 102
rect 190 98 194 102
rect 158 78 162 82
rect 126 68 130 72
rect 86 58 90 62
rect 214 118 218 122
rect 230 108 234 112
rect 222 78 226 82
rect 246 68 250 72
rect 430 818 434 822
rect 446 838 450 842
rect 462 838 466 842
rect 438 778 442 782
rect 454 748 458 752
rect 438 718 442 722
rect 422 668 426 672
rect 518 898 522 902
rect 518 888 522 892
rect 566 1048 570 1052
rect 614 1058 618 1062
rect 638 1058 642 1062
rect 654 1058 658 1062
rect 606 1048 610 1052
rect 646 1048 650 1052
rect 614 1008 618 1012
rect 646 1038 650 1042
rect 630 1028 634 1032
rect 678 1018 682 1022
rect 622 968 626 972
rect 646 968 650 972
rect 630 948 634 952
rect 702 948 706 952
rect 558 938 562 942
rect 582 928 586 932
rect 550 918 554 922
rect 598 918 602 922
rect 534 888 538 892
rect 646 908 650 912
rect 598 898 602 902
rect 590 888 594 892
rect 702 898 706 902
rect 622 888 626 892
rect 566 878 570 882
rect 694 878 698 882
rect 878 1318 882 1322
rect 894 1318 898 1322
rect 814 1308 818 1312
rect 838 1308 842 1312
rect 890 1303 894 1307
rect 897 1303 901 1307
rect 854 1278 858 1282
rect 862 1268 866 1272
rect 750 1148 754 1152
rect 782 1148 786 1152
rect 758 1128 762 1132
rect 774 1068 778 1072
rect 734 998 738 1002
rect 830 1168 834 1172
rect 958 1388 962 1392
rect 958 1338 962 1342
rect 1094 1558 1098 1562
rect 1118 1548 1122 1552
rect 1182 1548 1186 1552
rect 1086 1488 1090 1492
rect 1070 1478 1074 1482
rect 1142 1538 1146 1542
rect 1134 1488 1138 1492
rect 1102 1468 1106 1472
rect 1150 1508 1154 1512
rect 1158 1498 1162 1502
rect 1550 1698 1554 1702
rect 1438 1688 1442 1692
rect 1566 1678 1570 1682
rect 1766 1678 1770 1682
rect 1502 1668 1506 1672
rect 1750 1668 1754 1672
rect 1326 1658 1330 1662
rect 1366 1658 1370 1662
rect 1422 1658 1426 1662
rect 1358 1648 1362 1652
rect 1278 1578 1282 1582
rect 1302 1578 1306 1582
rect 1334 1548 1338 1552
rect 1238 1528 1242 1532
rect 1270 1528 1274 1532
rect 1190 1468 1194 1472
rect 1246 1468 1250 1472
rect 1126 1458 1130 1462
rect 1038 1388 1042 1392
rect 1030 1368 1034 1372
rect 1070 1378 1074 1382
rect 1078 1358 1082 1362
rect 1174 1438 1178 1442
rect 1150 1378 1154 1382
rect 1046 1348 1050 1352
rect 1070 1348 1074 1352
rect 1142 1348 1146 1352
rect 1022 1338 1026 1342
rect 1014 1328 1018 1332
rect 926 1158 930 1162
rect 846 1148 850 1152
rect 910 1148 914 1152
rect 1038 1298 1042 1302
rect 1086 1328 1090 1332
rect 1078 1298 1082 1302
rect 1102 1298 1106 1302
rect 1070 1288 1074 1292
rect 966 1278 970 1282
rect 1062 1278 1066 1282
rect 958 1268 962 1272
rect 1022 1268 1026 1272
rect 1270 1448 1274 1452
rect 1206 1418 1210 1422
rect 1286 1538 1290 1542
rect 1350 1518 1354 1522
rect 1294 1508 1298 1512
rect 1386 1603 1390 1607
rect 1393 1603 1397 1607
rect 1398 1558 1402 1562
rect 1478 1548 1482 1552
rect 1462 1538 1466 1542
rect 1422 1528 1426 1532
rect 1310 1478 1314 1482
rect 1342 1468 1346 1472
rect 1398 1478 1402 1482
rect 1310 1458 1314 1462
rect 1326 1458 1330 1462
rect 1358 1458 1362 1462
rect 1278 1388 1282 1392
rect 1326 1368 1330 1372
rect 1342 1358 1346 1362
rect 1270 1348 1274 1352
rect 1302 1348 1306 1352
rect 1158 1338 1162 1342
rect 1198 1338 1202 1342
rect 1286 1338 1290 1342
rect 1190 1328 1194 1332
rect 1238 1328 1242 1332
rect 1150 1308 1154 1312
rect 1166 1288 1170 1292
rect 1294 1308 1298 1312
rect 1270 1288 1274 1292
rect 1158 1278 1162 1282
rect 1206 1268 1210 1272
rect 1238 1268 1242 1272
rect 1278 1268 1282 1272
rect 998 1258 1002 1262
rect 1030 1258 1034 1262
rect 1062 1258 1066 1262
rect 1386 1403 1390 1407
rect 1393 1403 1397 1407
rect 1318 1328 1322 1332
rect 1350 1328 1354 1332
rect 1310 1298 1314 1302
rect 1310 1278 1314 1282
rect 1318 1268 1322 1272
rect 1342 1268 1346 1272
rect 1358 1268 1362 1272
rect 966 1208 970 1212
rect 958 1188 962 1192
rect 974 1178 978 1182
rect 942 1168 946 1172
rect 958 1168 962 1172
rect 966 1168 970 1172
rect 862 1138 866 1142
rect 830 1128 834 1132
rect 814 1118 818 1122
rect 806 1098 810 1102
rect 934 1128 938 1132
rect 878 1118 882 1122
rect 890 1103 894 1107
rect 897 1103 901 1107
rect 822 1068 826 1072
rect 862 1068 866 1072
rect 790 1028 794 1032
rect 766 968 770 972
rect 734 958 738 962
rect 734 938 738 942
rect 742 918 746 922
rect 758 918 762 922
rect 750 898 754 902
rect 566 868 570 872
rect 662 868 666 872
rect 686 868 690 872
rect 526 848 530 852
rect 534 798 538 802
rect 518 778 522 782
rect 502 758 506 762
rect 502 748 506 752
rect 486 688 490 692
rect 574 858 578 862
rect 622 858 626 862
rect 678 858 682 862
rect 702 858 706 862
rect 566 828 570 832
rect 558 768 562 772
rect 550 758 554 762
rect 614 758 618 762
rect 574 738 578 742
rect 542 718 546 722
rect 598 718 602 722
rect 574 708 578 712
rect 558 698 562 702
rect 486 678 490 682
rect 534 678 538 682
rect 454 668 458 672
rect 510 668 514 672
rect 430 658 434 662
rect 550 668 554 672
rect 494 658 498 662
rect 566 638 570 642
rect 438 628 442 632
rect 478 628 482 632
rect 370 603 374 607
rect 377 603 381 607
rect 334 558 338 562
rect 406 548 410 552
rect 318 528 322 532
rect 350 488 354 492
rect 270 478 274 482
rect 526 598 530 602
rect 446 578 450 582
rect 462 568 466 572
rect 502 558 506 562
rect 558 558 562 562
rect 470 548 474 552
rect 414 498 418 502
rect 278 468 282 472
rect 382 468 386 472
rect 318 458 322 462
rect 358 438 362 442
rect 286 418 290 422
rect 286 368 290 372
rect 342 368 346 372
rect 286 358 290 362
rect 302 338 306 342
rect 350 358 354 362
rect 370 403 374 407
rect 377 403 381 407
rect 406 358 410 362
rect 294 328 298 332
rect 366 328 370 332
rect 286 288 290 292
rect 310 288 314 292
rect 374 288 378 292
rect 422 338 426 342
rect 446 508 450 512
rect 494 548 498 552
rect 518 548 522 552
rect 542 548 546 552
rect 566 548 570 552
rect 486 528 490 532
rect 502 528 506 532
rect 510 528 514 532
rect 454 498 458 502
rect 438 488 442 492
rect 454 478 458 482
rect 454 408 458 412
rect 446 398 450 402
rect 558 518 562 522
rect 534 498 538 502
rect 526 468 530 472
rect 550 468 554 472
rect 462 368 466 372
rect 486 368 490 372
rect 510 368 514 372
rect 438 318 442 322
rect 470 338 474 342
rect 502 338 506 342
rect 494 328 498 332
rect 430 278 434 282
rect 430 268 434 272
rect 454 268 458 272
rect 406 258 410 262
rect 342 218 346 222
rect 374 218 378 222
rect 318 138 322 142
rect 278 88 282 92
rect 370 203 374 207
rect 377 203 381 207
rect 422 248 426 252
rect 374 188 378 192
rect 414 188 418 192
rect 390 148 394 152
rect 414 148 418 152
rect 462 248 466 252
rect 486 258 490 262
rect 542 368 546 372
rect 550 368 554 372
rect 550 358 554 362
rect 526 328 530 332
rect 534 328 538 332
rect 534 318 538 322
rect 550 288 554 292
rect 510 258 514 262
rect 550 258 554 262
rect 558 258 562 262
rect 494 228 498 232
rect 502 228 506 232
rect 502 218 506 222
rect 510 218 514 222
rect 518 218 522 222
rect 414 138 418 142
rect 374 128 378 132
rect 446 128 450 132
rect 510 148 514 152
rect 646 848 650 852
rect 646 838 650 842
rect 694 838 698 842
rect 662 818 666 822
rect 694 818 698 822
rect 718 818 722 822
rect 630 778 634 782
rect 662 758 666 762
rect 638 748 642 752
rect 630 728 634 732
rect 646 698 650 702
rect 622 668 626 672
rect 638 668 642 672
rect 726 798 730 802
rect 830 1018 834 1022
rect 862 998 866 1002
rect 910 988 914 992
rect 878 978 882 982
rect 814 968 818 972
rect 806 938 810 942
rect 774 858 778 862
rect 766 838 770 842
rect 742 818 746 822
rect 758 808 762 812
rect 734 778 738 782
rect 742 778 746 782
rect 734 768 738 772
rect 694 748 698 752
rect 750 748 754 752
rect 678 738 682 742
rect 702 728 706 732
rect 726 698 730 702
rect 806 838 810 842
rect 918 948 922 952
rect 830 928 834 932
rect 830 888 834 892
rect 838 888 842 892
rect 890 903 894 907
rect 897 903 901 907
rect 846 868 850 872
rect 782 788 786 792
rect 830 858 834 862
rect 942 988 946 992
rect 926 938 930 942
rect 830 778 834 782
rect 782 718 786 722
rect 774 708 778 712
rect 670 678 674 682
rect 662 658 666 662
rect 678 658 682 662
rect 598 648 602 652
rect 606 638 610 642
rect 582 558 586 562
rect 598 488 602 492
rect 670 588 674 592
rect 622 558 626 562
rect 614 528 618 532
rect 622 518 626 522
rect 646 518 650 522
rect 614 478 618 482
rect 654 468 658 472
rect 678 538 682 542
rect 742 658 746 662
rect 718 618 722 622
rect 798 688 802 692
rect 774 598 778 602
rect 734 558 738 562
rect 782 548 786 552
rect 702 538 706 542
rect 670 528 674 532
rect 694 528 698 532
rect 734 528 738 532
rect 686 488 690 492
rect 686 468 690 472
rect 598 458 602 462
rect 630 458 634 462
rect 574 438 578 442
rect 654 378 658 382
rect 670 368 674 372
rect 646 358 650 362
rect 654 358 658 362
rect 678 358 682 362
rect 582 348 586 352
rect 630 338 634 342
rect 638 338 642 342
rect 598 328 602 332
rect 590 298 594 302
rect 718 478 722 482
rect 718 448 722 452
rect 710 368 714 372
rect 702 358 706 362
rect 686 348 690 352
rect 694 338 698 342
rect 686 328 690 332
rect 638 318 642 322
rect 630 298 634 302
rect 598 278 602 282
rect 622 278 626 282
rect 614 268 618 272
rect 654 298 658 302
rect 694 318 698 322
rect 646 288 650 292
rect 678 288 682 292
rect 598 258 602 262
rect 614 258 618 262
rect 622 258 626 262
rect 630 258 634 262
rect 638 258 642 262
rect 606 238 610 242
rect 614 228 618 232
rect 606 158 610 162
rect 494 138 498 142
rect 334 88 338 92
rect 494 88 498 92
rect 374 78 378 82
rect 414 78 418 82
rect 278 68 282 72
rect 294 68 298 72
rect 206 58 210 62
rect 238 58 242 62
rect 262 58 266 62
rect 526 138 530 142
rect 558 138 562 142
rect 574 138 578 142
rect 590 138 594 142
rect 598 128 602 132
rect 526 78 530 82
rect 470 58 474 62
rect 502 58 506 62
rect 558 58 562 62
rect 198 48 202 52
rect 566 8 570 12
rect 370 3 374 7
rect 377 3 381 7
rect 726 358 730 362
rect 718 348 722 352
rect 710 278 714 282
rect 702 268 706 272
rect 678 248 682 252
rect 670 168 674 172
rect 686 218 690 222
rect 686 158 690 162
rect 654 148 658 152
rect 662 88 666 92
rect 694 88 698 92
rect 630 58 634 62
rect 630 8 634 12
rect 646 8 650 12
rect 758 528 762 532
rect 750 368 754 372
rect 766 468 770 472
rect 790 518 794 522
rect 870 838 874 842
rect 846 748 850 752
rect 822 738 826 742
rect 814 718 818 722
rect 814 658 818 662
rect 854 718 858 722
rect 846 708 850 712
rect 910 788 914 792
rect 918 758 922 762
rect 1006 1248 1010 1252
rect 1038 1248 1042 1252
rect 1022 1238 1026 1242
rect 990 1228 994 1232
rect 990 1168 994 1172
rect 982 1138 986 1142
rect 966 1128 970 1132
rect 1014 1118 1018 1122
rect 990 1108 994 1112
rect 990 1098 994 1102
rect 974 1078 978 1082
rect 982 1078 986 1082
rect 1142 1238 1146 1242
rect 1126 1168 1130 1172
rect 1406 1318 1410 1322
rect 1454 1518 1458 1522
rect 1558 1588 1562 1592
rect 1526 1518 1530 1522
rect 1470 1478 1474 1482
rect 1598 1658 1602 1662
rect 1670 1658 1674 1662
rect 1726 1658 1730 1662
rect 1702 1648 1706 1652
rect 1686 1638 1690 1642
rect 1646 1608 1650 1612
rect 1654 1608 1658 1612
rect 1574 1558 1578 1562
rect 1566 1518 1570 1522
rect 1558 1498 1562 1502
rect 1582 1538 1586 1542
rect 1622 1528 1626 1532
rect 1710 1558 1714 1562
rect 1726 1558 1730 1562
rect 1638 1518 1642 1522
rect 1678 1518 1682 1522
rect 1614 1508 1618 1512
rect 1574 1488 1578 1492
rect 1718 1508 1722 1512
rect 1734 1498 1738 1502
rect 1646 1488 1650 1492
rect 1702 1488 1706 1492
rect 1550 1478 1554 1482
rect 1638 1478 1642 1482
rect 1526 1468 1530 1472
rect 1542 1468 1546 1472
rect 1566 1468 1570 1472
rect 1446 1448 1450 1452
rect 1438 1348 1442 1352
rect 1486 1448 1490 1452
rect 1550 1458 1554 1462
rect 1598 1458 1602 1462
rect 1686 1458 1690 1462
rect 1566 1448 1570 1452
rect 1494 1428 1498 1432
rect 1486 1378 1490 1382
rect 1470 1338 1474 1342
rect 1534 1338 1538 1342
rect 1430 1328 1434 1332
rect 1478 1308 1482 1312
rect 1510 1308 1514 1312
rect 1510 1288 1514 1292
rect 1518 1288 1522 1292
rect 1502 1278 1506 1282
rect 1470 1268 1474 1272
rect 1630 1448 1634 1452
rect 1766 1658 1770 1662
rect 1798 1658 1802 1662
rect 1790 1578 1794 1582
rect 1790 1568 1794 1572
rect 1750 1478 1754 1482
rect 1702 1418 1706 1422
rect 1742 1418 1746 1422
rect 1598 1378 1602 1382
rect 1638 1378 1642 1382
rect 1566 1368 1570 1372
rect 1686 1368 1690 1372
rect 1598 1358 1602 1362
rect 1630 1358 1634 1362
rect 1662 1358 1666 1362
rect 1574 1338 1578 1342
rect 1542 1328 1546 1332
rect 1598 1318 1602 1322
rect 1606 1298 1610 1302
rect 1374 1258 1378 1262
rect 1358 1248 1362 1252
rect 1334 1238 1338 1242
rect 1286 1228 1290 1232
rect 1294 1228 1298 1232
rect 1334 1228 1338 1232
rect 1214 1158 1218 1162
rect 1326 1158 1330 1162
rect 1046 1148 1050 1152
rect 998 1058 1002 1062
rect 1030 1058 1034 1062
rect 1006 1038 1010 1042
rect 966 1018 970 1022
rect 998 988 1002 992
rect 998 968 1002 972
rect 958 958 962 962
rect 966 958 970 962
rect 966 938 970 942
rect 958 928 962 932
rect 950 868 954 872
rect 982 928 986 932
rect 998 918 1002 922
rect 998 898 1002 902
rect 1046 968 1050 972
rect 1078 1128 1082 1132
rect 1094 1118 1098 1122
rect 1070 1108 1074 1112
rect 1094 1088 1098 1092
rect 1102 1088 1106 1092
rect 1070 1068 1074 1072
rect 1126 1058 1130 1062
rect 1150 1138 1154 1142
rect 1326 1138 1330 1142
rect 1214 1128 1218 1132
rect 1150 1118 1154 1122
rect 1262 1068 1266 1072
rect 1158 1058 1162 1062
rect 1310 1058 1314 1062
rect 1206 1038 1210 1042
rect 1230 1038 1234 1042
rect 1142 988 1146 992
rect 1062 948 1066 952
rect 1126 948 1130 952
rect 1046 938 1050 942
rect 1022 878 1026 882
rect 990 868 994 872
rect 1014 868 1018 872
rect 958 858 962 862
rect 974 858 978 862
rect 990 858 994 862
rect 1030 858 1034 862
rect 950 848 954 852
rect 934 838 938 842
rect 966 838 970 842
rect 974 778 978 782
rect 1006 818 1010 822
rect 1006 798 1010 802
rect 1022 788 1026 792
rect 1006 768 1010 772
rect 998 748 1002 752
rect 966 738 970 742
rect 974 738 978 742
rect 890 703 894 707
rect 897 703 901 707
rect 950 708 954 712
rect 926 688 930 692
rect 910 678 914 682
rect 854 668 858 672
rect 854 648 858 652
rect 862 648 866 652
rect 846 638 850 642
rect 918 648 922 652
rect 894 618 898 622
rect 838 608 842 612
rect 854 608 858 612
rect 838 598 842 602
rect 918 558 922 562
rect 814 538 818 542
rect 806 518 810 522
rect 814 458 818 462
rect 814 448 818 452
rect 814 428 818 432
rect 782 418 786 422
rect 774 348 778 352
rect 758 328 762 332
rect 758 318 762 322
rect 750 268 754 272
rect 766 268 770 272
rect 742 258 746 262
rect 750 238 754 242
rect 750 198 754 202
rect 806 388 810 392
rect 790 378 794 382
rect 902 528 906 532
rect 878 518 882 522
rect 838 468 842 472
rect 890 503 894 507
rect 897 503 901 507
rect 910 488 914 492
rect 1006 728 1010 732
rect 1022 728 1026 732
rect 998 708 1002 712
rect 1062 868 1066 872
rect 1150 938 1154 942
rect 1174 928 1178 932
rect 1158 918 1162 922
rect 1222 948 1226 952
rect 1286 1018 1290 1022
rect 1358 1138 1362 1142
rect 1358 1128 1362 1132
rect 1342 1078 1346 1082
rect 1406 1218 1410 1222
rect 1386 1203 1390 1207
rect 1393 1203 1397 1207
rect 1398 1168 1402 1172
rect 1462 1138 1466 1142
rect 1438 1128 1442 1132
rect 1446 1128 1450 1132
rect 1526 1128 1530 1132
rect 1550 1128 1554 1132
rect 1374 1118 1378 1122
rect 1438 1078 1442 1082
rect 1430 1068 1434 1072
rect 1438 1048 1442 1052
rect 1350 1028 1354 1032
rect 1334 1008 1338 1012
rect 1334 988 1338 992
rect 1326 958 1330 962
rect 1238 908 1242 912
rect 1278 918 1282 922
rect 1386 1003 1390 1007
rect 1393 1003 1397 1007
rect 1374 958 1378 962
rect 1374 938 1378 942
rect 1358 918 1362 922
rect 1470 1118 1474 1122
rect 1510 1118 1514 1122
rect 1462 1068 1466 1072
rect 1478 1068 1482 1072
rect 1494 1068 1498 1072
rect 1486 1058 1490 1062
rect 1470 1008 1474 1012
rect 1486 958 1490 962
rect 1430 918 1434 922
rect 1406 908 1410 912
rect 1630 1278 1634 1282
rect 1670 1348 1674 1352
rect 1670 1328 1674 1332
rect 1678 1328 1682 1332
rect 1646 1278 1650 1282
rect 1670 1278 1674 1282
rect 1638 1268 1642 1272
rect 1654 1258 1658 1262
rect 1662 1258 1666 1262
rect 1622 1248 1626 1252
rect 1598 1238 1602 1242
rect 1622 1208 1626 1212
rect 1614 1178 1618 1182
rect 1598 1158 1602 1162
rect 1606 1148 1610 1152
rect 1614 1138 1618 1142
rect 1574 1098 1578 1102
rect 1550 1058 1554 1062
rect 1534 958 1538 962
rect 1526 908 1530 912
rect 1510 898 1514 902
rect 1478 888 1482 892
rect 1446 878 1450 882
rect 1494 868 1498 872
rect 1670 1208 1674 1212
rect 1670 1178 1674 1182
rect 1654 1158 1658 1162
rect 1630 1138 1634 1142
rect 1638 1128 1642 1132
rect 1646 1128 1650 1132
rect 1622 1098 1626 1102
rect 1622 1088 1626 1092
rect 1686 1268 1690 1272
rect 1742 1408 1746 1412
rect 1734 1388 1738 1392
rect 1726 1338 1730 1342
rect 1710 1318 1714 1322
rect 1734 1278 1738 1282
rect 1758 1368 1762 1372
rect 1758 1358 1762 1362
rect 1774 1508 1778 1512
rect 1774 1418 1778 1422
rect 1782 1348 1786 1352
rect 1782 1328 1786 1332
rect 1766 1278 1770 1282
rect 1718 1258 1722 1262
rect 1694 1178 1698 1182
rect 1710 1168 1714 1172
rect 1734 1248 1738 1252
rect 1750 1218 1754 1222
rect 1694 1148 1698 1152
rect 1702 1138 1706 1142
rect 1686 1088 1690 1092
rect 1630 1068 1634 1072
rect 1638 1068 1642 1072
rect 1646 1068 1650 1072
rect 1662 1068 1666 1072
rect 1686 1068 1690 1072
rect 1702 1068 1706 1072
rect 1622 1058 1626 1062
rect 1598 1048 1602 1052
rect 1630 1018 1634 1022
rect 1630 1008 1634 1012
rect 1590 998 1594 1002
rect 1598 988 1602 992
rect 1606 968 1610 972
rect 1654 1048 1658 1052
rect 1654 1018 1658 1022
rect 1638 948 1642 952
rect 1582 938 1586 942
rect 1622 938 1626 942
rect 1646 918 1650 922
rect 1614 888 1618 892
rect 1630 888 1634 892
rect 1582 878 1586 882
rect 1638 878 1642 882
rect 1590 868 1594 872
rect 1638 868 1642 872
rect 1670 1048 1674 1052
rect 1662 918 1666 922
rect 1670 888 1674 892
rect 1694 1058 1698 1062
rect 1710 958 1714 962
rect 1710 878 1714 882
rect 1166 858 1170 862
rect 1230 858 1234 862
rect 1254 858 1258 862
rect 1158 848 1162 852
rect 1174 848 1178 852
rect 1190 848 1194 852
rect 1142 838 1146 842
rect 1230 848 1234 852
rect 1206 808 1210 812
rect 1110 788 1114 792
rect 1142 788 1146 792
rect 1054 778 1058 782
rect 1086 778 1090 782
rect 1142 778 1146 782
rect 1134 768 1138 772
rect 1182 768 1186 772
rect 1070 748 1074 752
rect 1038 708 1042 712
rect 982 688 986 692
rect 998 688 1002 692
rect 1014 688 1018 692
rect 982 668 986 672
rect 982 598 986 602
rect 942 548 946 552
rect 974 548 978 552
rect 966 538 970 542
rect 1014 668 1018 672
rect 1038 668 1042 672
rect 1038 628 1042 632
rect 1006 598 1010 602
rect 1006 578 1010 582
rect 990 548 994 552
rect 974 528 978 532
rect 974 488 978 492
rect 926 478 930 482
rect 982 478 986 482
rect 998 538 1002 542
rect 1030 508 1034 512
rect 934 468 938 472
rect 974 458 978 462
rect 894 438 898 442
rect 830 358 834 362
rect 838 358 842 362
rect 822 348 826 352
rect 798 328 802 332
rect 814 328 818 332
rect 798 288 802 292
rect 830 288 834 292
rect 806 278 810 282
rect 798 268 802 272
rect 806 188 810 192
rect 790 158 794 162
rect 750 148 754 152
rect 718 138 722 142
rect 734 138 738 142
rect 718 68 722 72
rect 782 78 786 82
rect 734 58 738 62
rect 774 58 778 62
rect 774 8 778 12
rect 790 8 794 12
rect 886 368 890 372
rect 918 368 922 372
rect 910 348 914 352
rect 878 338 882 342
rect 870 328 874 332
rect 854 318 858 322
rect 890 303 894 307
rect 897 303 901 307
rect 942 388 946 392
rect 990 388 994 392
rect 974 358 978 362
rect 958 348 962 352
rect 918 288 922 292
rect 926 288 930 292
rect 886 268 890 272
rect 958 268 962 272
rect 1014 478 1018 482
rect 1062 738 1066 742
rect 1102 718 1106 722
rect 1102 698 1106 702
rect 1078 688 1082 692
rect 1110 688 1114 692
rect 1190 718 1194 722
rect 1182 708 1186 712
rect 1070 668 1074 672
rect 1166 678 1170 682
rect 1174 668 1178 672
rect 1054 648 1058 652
rect 1158 648 1162 652
rect 1062 638 1066 642
rect 1102 598 1106 602
rect 1062 547 1066 551
rect 1150 568 1154 572
rect 1222 778 1226 782
rect 1238 778 1242 782
rect 1238 768 1242 772
rect 1246 768 1250 772
rect 1318 818 1322 822
rect 1326 818 1330 822
rect 1278 808 1282 812
rect 1286 768 1290 772
rect 1310 768 1314 772
rect 1270 748 1274 752
rect 1294 748 1298 752
rect 1238 708 1242 712
rect 1214 678 1218 682
rect 1214 668 1218 672
rect 1238 668 1242 672
rect 1182 658 1186 662
rect 1230 658 1234 662
rect 1198 648 1202 652
rect 1182 588 1186 592
rect 1118 548 1122 552
rect 1142 548 1146 552
rect 1190 578 1194 582
rect 1214 618 1218 622
rect 1238 598 1242 602
rect 1190 548 1194 552
rect 1206 548 1210 552
rect 1054 518 1058 522
rect 1102 518 1106 522
rect 1078 498 1082 502
rect 1094 488 1098 492
rect 1046 478 1050 482
rect 1086 478 1090 482
rect 1030 458 1034 462
rect 1006 428 1010 432
rect 1046 428 1050 432
rect 1014 398 1018 402
rect 1030 388 1034 392
rect 1046 368 1050 372
rect 1006 358 1010 362
rect 1038 328 1042 332
rect 1006 288 1010 292
rect 1062 378 1066 382
rect 1070 348 1074 352
rect 1166 508 1170 512
rect 1182 498 1186 502
rect 1238 538 1242 542
rect 1222 498 1226 502
rect 1214 488 1218 492
rect 1206 478 1210 482
rect 1126 468 1130 472
rect 1238 488 1242 492
rect 1222 458 1226 462
rect 1238 458 1242 462
rect 1166 448 1170 452
rect 1182 448 1186 452
rect 1206 448 1210 452
rect 1094 368 1098 372
rect 1062 338 1066 342
rect 1086 338 1090 342
rect 1078 318 1082 322
rect 1078 308 1082 312
rect 974 258 978 262
rect 1038 258 1042 262
rect 966 208 970 212
rect 998 208 1002 212
rect 910 188 914 192
rect 878 168 882 172
rect 862 158 866 162
rect 958 158 962 162
rect 982 188 986 192
rect 1070 188 1074 192
rect 1006 168 1010 172
rect 1038 158 1042 162
rect 926 148 930 152
rect 950 148 954 152
rect 890 103 894 107
rect 897 103 901 107
rect 1142 328 1146 332
rect 1270 698 1274 702
rect 1270 648 1274 652
rect 1310 608 1314 612
rect 1302 548 1306 552
rect 1278 518 1282 522
rect 1278 468 1282 472
rect 1334 808 1338 812
rect 1326 758 1330 762
rect 1326 728 1330 732
rect 1374 848 1378 852
rect 1386 803 1390 807
rect 1393 803 1397 807
rect 1358 798 1362 802
rect 1350 758 1354 762
rect 1390 778 1394 782
rect 1374 768 1378 772
rect 1342 718 1346 722
rect 1358 678 1362 682
rect 1342 668 1346 672
rect 1350 658 1354 662
rect 1358 658 1362 662
rect 1382 708 1386 712
rect 1422 748 1426 752
rect 1430 748 1434 752
rect 1414 688 1418 692
rect 1414 668 1418 672
rect 1446 728 1450 732
rect 1470 718 1474 722
rect 1438 678 1442 682
rect 1374 628 1378 632
rect 1366 598 1370 602
rect 1326 578 1330 582
rect 1334 558 1338 562
rect 1350 548 1354 552
rect 1366 518 1370 522
rect 1366 478 1370 482
rect 1310 468 1314 472
rect 1334 468 1338 472
rect 1342 468 1346 472
rect 1270 458 1274 462
rect 1198 348 1202 352
rect 1222 348 1226 352
rect 1206 338 1210 342
rect 1222 328 1226 332
rect 1238 308 1242 312
rect 1254 308 1258 312
rect 1270 338 1274 342
rect 1190 288 1194 292
rect 1110 258 1114 262
rect 1142 258 1146 262
rect 1158 258 1162 262
rect 1166 248 1170 252
rect 1126 208 1130 212
rect 1118 198 1122 202
rect 1102 168 1106 172
rect 1246 278 1250 282
rect 1262 278 1266 282
rect 1214 268 1218 272
rect 1326 448 1330 452
rect 1366 438 1370 442
rect 1326 408 1330 412
rect 1342 328 1346 332
rect 1386 603 1390 607
rect 1393 603 1397 607
rect 1430 648 1434 652
rect 1430 618 1434 622
rect 1446 618 1450 622
rect 1422 578 1426 582
rect 1390 558 1394 562
rect 1430 558 1434 562
rect 1438 558 1442 562
rect 1382 548 1386 552
rect 1414 548 1418 552
rect 1422 538 1426 542
rect 1558 718 1562 722
rect 1550 698 1554 702
rect 1542 688 1546 692
rect 1478 648 1482 652
rect 1462 638 1466 642
rect 1526 648 1530 652
rect 1550 648 1554 652
rect 1542 628 1546 632
rect 1518 598 1522 602
rect 1478 578 1482 582
rect 1494 568 1498 572
rect 1454 528 1458 532
rect 1438 508 1442 512
rect 1462 478 1466 482
rect 1386 403 1390 407
rect 1393 403 1397 407
rect 1574 588 1578 592
rect 1574 568 1578 572
rect 1558 548 1562 552
rect 1558 538 1562 542
rect 1542 518 1546 522
rect 1534 508 1538 512
rect 1550 508 1554 512
rect 1502 458 1506 462
rect 1478 448 1482 452
rect 1486 418 1490 422
rect 1406 388 1410 392
rect 1414 388 1418 392
rect 1374 318 1378 322
rect 1390 318 1394 322
rect 1302 288 1306 292
rect 1430 308 1434 312
rect 1326 268 1330 272
rect 1270 258 1274 262
rect 1182 208 1186 212
rect 1142 158 1146 162
rect 1158 158 1162 162
rect 1174 158 1178 162
rect 1094 148 1098 152
rect 1174 148 1178 152
rect 1238 248 1242 252
rect 1214 208 1218 212
rect 1222 158 1226 162
rect 1206 148 1210 152
rect 1238 148 1242 152
rect 1302 248 1306 252
rect 1366 238 1370 242
rect 1374 228 1378 232
rect 1366 218 1370 222
rect 1366 168 1370 172
rect 1302 148 1306 152
rect 1150 138 1154 142
rect 1174 128 1178 132
rect 1190 128 1194 132
rect 1126 118 1130 122
rect 966 98 970 102
rect 1046 88 1050 92
rect 1118 88 1122 92
rect 830 68 834 72
rect 902 68 906 72
rect 862 58 866 62
rect 934 58 938 62
rect 894 48 898 52
rect 1022 59 1026 63
rect 1134 98 1138 102
rect 1238 118 1242 122
rect 1230 108 1234 112
rect 1270 88 1274 92
rect 1198 78 1202 82
rect 1214 78 1218 82
rect 1230 78 1234 82
rect 1166 58 1170 62
rect 1078 38 1082 42
rect 942 8 946 12
rect 958 8 962 12
rect 1222 58 1226 62
rect 1294 78 1298 82
rect 1358 78 1362 82
rect 1386 203 1390 207
rect 1393 203 1397 207
rect 1414 228 1418 232
rect 1406 178 1410 182
rect 1406 168 1410 172
rect 1438 288 1442 292
rect 1446 288 1450 292
rect 1470 318 1474 322
rect 1462 248 1466 252
rect 1454 218 1458 222
rect 1518 398 1522 402
rect 1542 448 1546 452
rect 1534 318 1538 322
rect 1566 508 1570 512
rect 1566 498 1570 502
rect 1558 438 1562 442
rect 1622 848 1626 852
rect 1622 748 1626 752
rect 1638 708 1642 712
rect 1638 688 1642 692
rect 1630 678 1634 682
rect 1670 838 1674 842
rect 1654 758 1658 762
rect 1662 738 1666 742
rect 1670 688 1674 692
rect 1686 858 1690 862
rect 1702 858 1706 862
rect 1734 1128 1738 1132
rect 1742 1108 1746 1112
rect 1758 1058 1762 1062
rect 1766 1048 1770 1052
rect 1798 1238 1802 1242
rect 1798 1208 1802 1212
rect 1798 1038 1802 1042
rect 1750 928 1754 932
rect 1734 918 1738 922
rect 1774 908 1778 912
rect 1726 878 1730 882
rect 1798 878 1802 882
rect 1782 868 1786 872
rect 1702 848 1706 852
rect 1718 848 1722 852
rect 1710 788 1714 792
rect 1686 748 1690 752
rect 1750 748 1754 752
rect 1686 718 1690 722
rect 1678 668 1682 672
rect 1606 658 1610 662
rect 1646 658 1650 662
rect 1598 638 1602 642
rect 1614 598 1618 602
rect 1598 578 1602 582
rect 1614 538 1618 542
rect 1614 508 1618 512
rect 1598 478 1602 482
rect 1598 468 1602 472
rect 1582 438 1586 442
rect 1630 638 1634 642
rect 1638 598 1642 602
rect 1654 558 1658 562
rect 1678 658 1682 662
rect 1726 658 1730 662
rect 1670 648 1674 652
rect 1702 618 1706 622
rect 1694 608 1698 612
rect 1686 568 1690 572
rect 1686 538 1690 542
rect 1710 588 1714 592
rect 1702 558 1706 562
rect 1662 488 1666 492
rect 1790 578 1794 582
rect 1662 478 1666 482
rect 1686 468 1690 472
rect 1622 418 1626 422
rect 1630 408 1634 412
rect 1646 408 1650 412
rect 1582 398 1586 402
rect 1614 348 1618 352
rect 1590 318 1594 322
rect 1534 268 1538 272
rect 1502 258 1506 262
rect 1582 258 1586 262
rect 1510 248 1514 252
rect 1566 228 1570 232
rect 1526 178 1530 182
rect 1470 168 1474 172
rect 1486 168 1490 172
rect 1486 158 1490 162
rect 1558 158 1562 162
rect 1382 148 1386 152
rect 1430 148 1434 152
rect 1518 148 1522 152
rect 1614 258 1618 262
rect 1598 188 1602 192
rect 1590 178 1594 182
rect 1462 138 1466 142
rect 1478 138 1482 142
rect 1446 128 1450 132
rect 1382 88 1386 92
rect 1406 78 1410 82
rect 1494 128 1498 132
rect 1606 88 1610 92
rect 1622 198 1626 202
rect 1638 358 1642 362
rect 1766 538 1770 542
rect 1750 518 1754 522
rect 1694 458 1698 462
rect 1694 448 1698 452
rect 1742 448 1746 452
rect 1670 398 1674 402
rect 1718 418 1722 422
rect 1718 398 1722 402
rect 1702 348 1706 352
rect 1646 318 1650 322
rect 1702 338 1706 342
rect 1694 298 1698 302
rect 1710 328 1714 332
rect 1774 508 1778 512
rect 1758 458 1762 462
rect 1766 438 1770 442
rect 1758 358 1762 362
rect 1782 368 1786 372
rect 1694 278 1698 282
rect 1734 268 1738 272
rect 1798 288 1802 292
rect 1742 258 1746 262
rect 1790 258 1794 262
rect 1734 248 1738 252
rect 1686 238 1690 242
rect 1718 238 1722 242
rect 1694 228 1698 232
rect 1694 218 1698 222
rect 1742 228 1746 232
rect 1662 158 1666 162
rect 1702 158 1706 162
rect 1726 158 1730 162
rect 1646 148 1650 152
rect 1630 138 1634 142
rect 1638 108 1642 112
rect 1462 68 1466 72
rect 1494 68 1498 72
rect 1534 68 1538 72
rect 1438 58 1442 62
rect 1502 58 1506 62
rect 1782 218 1786 222
rect 1790 168 1794 172
rect 1758 158 1762 162
rect 1774 148 1778 152
rect 1702 128 1706 132
rect 1766 108 1770 112
rect 1694 98 1698 102
rect 1718 98 1722 102
rect 1790 98 1794 102
rect 1678 88 1682 92
rect 1710 78 1714 82
rect 1726 68 1730 72
rect 1470 48 1474 52
rect 1386 3 1390 7
rect 1393 3 1397 7
<< metal3 >>
rect 1830 1718 1834 1722
rect 1830 1711 1833 1718
rect 1822 1708 1833 1711
rect 888 1703 890 1707
rect 894 1703 897 1707
rect 902 1703 904 1707
rect 1822 1701 1825 1708
rect 1554 1698 1825 1701
rect 1830 1698 1834 1702
rect 18 1688 150 1691
rect 154 1688 318 1691
rect 434 1688 518 1691
rect 1830 1691 1833 1698
rect 1766 1688 1833 1691
rect 706 1678 718 1681
rect 818 1678 830 1681
rect 858 1678 870 1681
rect 1254 1681 1257 1688
rect 1438 1681 1441 1688
rect 1766 1682 1769 1688
rect 1254 1678 1566 1681
rect 1830 1678 1834 1682
rect 342 1671 345 1678
rect 342 1668 422 1671
rect 426 1668 494 1671
rect 1422 1668 1502 1671
rect 1830 1671 1833 1678
rect 1754 1668 1833 1671
rect 62 1662 65 1668
rect 66 1658 366 1661
rect 370 1658 406 1661
rect 494 1661 497 1668
rect 1422 1662 1425 1668
rect 418 1658 465 1661
rect 494 1658 542 1661
rect 546 1658 614 1661
rect 882 1658 1022 1661
rect 1026 1658 1038 1661
rect 1050 1658 1110 1661
rect 1330 1658 1366 1661
rect 1594 1658 1598 1661
rect 1650 1658 1670 1661
rect 1674 1658 1726 1661
rect 1762 1658 1766 1661
rect 1830 1661 1834 1662
rect 1802 1658 1834 1661
rect 38 1651 41 1658
rect 462 1652 465 1658
rect 38 1648 94 1651
rect 810 1648 918 1651
rect 922 1648 934 1651
rect 946 1648 1254 1651
rect 1362 1648 1702 1651
rect 386 1638 446 1641
rect 450 1638 878 1641
rect 1010 1638 1014 1641
rect 1690 1638 1742 1641
rect 1830 1641 1834 1642
rect 1786 1638 1834 1641
rect 346 1628 598 1631
rect 602 1628 742 1631
rect 746 1628 1318 1631
rect 154 1618 726 1621
rect 1646 1618 1694 1621
rect 1830 1621 1834 1622
rect 1802 1618 1834 1621
rect 1646 1612 1649 1618
rect 66 1608 126 1611
rect 130 1608 222 1611
rect 226 1608 286 1611
rect 368 1603 370 1607
rect 374 1603 377 1607
rect 382 1603 384 1607
rect 694 1602 697 1608
rect 1384 1603 1386 1607
rect 1390 1603 1393 1607
rect 1398 1603 1400 1607
rect 1654 1602 1657 1608
rect 1830 1601 1834 1602
rect 1794 1598 1834 1601
rect 266 1588 574 1591
rect 642 1588 934 1591
rect 1178 1588 1558 1591
rect 330 1578 542 1581
rect 730 1578 878 1581
rect 882 1578 1278 1581
rect 1282 1578 1302 1581
rect 1830 1581 1834 1582
rect 1794 1578 1834 1581
rect 1058 1568 1070 1571
rect 1130 1568 1142 1571
rect 1146 1568 1153 1571
rect 1794 1568 1798 1571
rect 194 1558 262 1561
rect 266 1558 598 1561
rect 602 1558 606 1561
rect 706 1558 806 1561
rect 1018 1558 1094 1561
rect 1682 1558 1710 1561
rect 1730 1558 1734 1561
rect 58 1548 206 1551
rect 210 1548 222 1551
rect 410 1548 598 1551
rect 702 1551 705 1558
rect 682 1548 705 1551
rect 794 1548 830 1551
rect 766 1542 769 1548
rect 874 1548 902 1551
rect 922 1548 1014 1551
rect 1122 1548 1182 1551
rect 1398 1551 1401 1558
rect 1338 1548 1401 1551
rect 1482 1548 1486 1551
rect 1574 1551 1577 1558
rect 1490 1548 1577 1551
rect 42 1538 126 1541
rect 154 1538 158 1541
rect 162 1538 190 1541
rect 482 1538 494 1541
rect 642 1538 726 1541
rect 1034 1538 1142 1541
rect 1146 1538 1286 1541
rect 1322 1538 1462 1541
rect 1586 1538 1625 1541
rect 114 1528 166 1531
rect 190 1531 193 1538
rect 1622 1532 1625 1538
rect 190 1528 518 1531
rect 738 1528 918 1531
rect 1010 1528 1238 1531
rect 1274 1528 1422 1531
rect 402 1518 502 1521
rect 698 1518 966 1521
rect 978 1518 1038 1521
rect 1050 1518 1350 1521
rect 1354 1518 1454 1521
rect 1530 1518 1566 1521
rect 1570 1518 1638 1521
rect 1682 1518 1726 1521
rect 514 1508 614 1511
rect 618 1508 734 1511
rect 1010 1508 1150 1511
rect 1154 1508 1294 1511
rect 1618 1508 1718 1511
rect 1722 1508 1774 1511
rect 888 1503 890 1507
rect 894 1503 897 1507
rect 902 1503 904 1507
rect 426 1498 430 1501
rect 434 1498 494 1501
rect 522 1498 806 1501
rect 810 1498 870 1501
rect 986 1498 1014 1501
rect 1026 1498 1158 1501
rect 1562 1498 1734 1501
rect 442 1488 566 1491
rect 570 1488 598 1491
rect 1090 1488 1134 1491
rect 1578 1488 1646 1491
rect 98 1478 110 1481
rect 114 1478 158 1481
rect 202 1478 622 1481
rect 990 1481 993 1488
rect 650 1478 993 1481
rect 1018 1478 1070 1481
rect 1314 1478 1398 1481
rect 1554 1478 1582 1481
rect 1702 1481 1705 1488
rect 1642 1478 1750 1481
rect 122 1468 134 1471
rect 138 1468 406 1471
rect 410 1468 422 1471
rect 426 1468 478 1471
rect 490 1468 494 1471
rect 626 1468 630 1471
rect 658 1468 662 1471
rect 858 1468 926 1471
rect 930 1468 934 1471
rect 938 1468 1030 1471
rect 1034 1468 1102 1471
rect 1106 1468 1190 1471
rect 1194 1468 1246 1471
rect 1470 1471 1473 1478
rect 1470 1468 1526 1471
rect 1546 1468 1558 1471
rect 1570 1468 1574 1471
rect 1342 1462 1345 1468
rect 1686 1462 1689 1468
rect 50 1458 126 1461
rect 258 1458 326 1461
rect 394 1458 526 1461
rect 546 1458 774 1461
rect 778 1458 822 1461
rect 826 1458 838 1461
rect 850 1458 934 1461
rect 1002 1458 1006 1461
rect 1042 1458 1126 1461
rect 1130 1458 1310 1461
rect 1346 1458 1358 1461
rect 1482 1458 1489 1461
rect 1554 1458 1598 1461
rect 194 1448 286 1451
rect 414 1448 422 1451
rect 426 1448 454 1451
rect 466 1448 606 1451
rect 610 1448 654 1451
rect 802 1448 814 1451
rect 818 1448 878 1451
rect 1174 1448 1270 1451
rect 1326 1451 1329 1458
rect 1486 1452 1489 1458
rect 1326 1448 1446 1451
rect 1570 1448 1630 1451
rect 462 1442 465 1448
rect 1174 1442 1177 1448
rect 178 1438 462 1441
rect 394 1428 422 1431
rect 810 1428 1494 1431
rect 686 1422 689 1428
rect 522 1418 606 1421
rect 794 1418 878 1421
rect 938 1418 1206 1421
rect 1706 1418 1742 1421
rect 1746 1418 1774 1421
rect 690 1408 694 1411
rect 1594 1408 1742 1411
rect 368 1403 370 1407
rect 374 1403 377 1407
rect 382 1403 384 1407
rect 1384 1403 1386 1407
rect 1390 1403 1393 1407
rect 1398 1403 1400 1407
rect 410 1388 598 1391
rect 602 1388 702 1391
rect 706 1388 774 1391
rect 962 1388 1038 1391
rect 1282 1388 1734 1391
rect 274 1378 366 1381
rect 658 1378 798 1381
rect 1002 1378 1070 1381
rect 1490 1378 1598 1381
rect 1602 1378 1638 1381
rect 1150 1372 1153 1378
rect 202 1368 254 1371
rect 266 1368 342 1371
rect 346 1368 558 1371
rect 562 1368 614 1371
rect 618 1368 646 1371
rect 1034 1368 1038 1371
rect 1330 1368 1566 1371
rect 1570 1368 1686 1371
rect 1754 1368 1758 1371
rect 154 1358 206 1361
rect 226 1358 230 1361
rect 282 1358 294 1361
rect 306 1358 310 1361
rect 578 1358 582 1361
rect 594 1358 598 1361
rect 662 1361 665 1368
rect 602 1358 665 1361
rect 722 1358 758 1361
rect 930 1358 1078 1361
rect 1602 1358 1630 1361
rect 1666 1358 1758 1361
rect 146 1348 230 1351
rect 242 1348 278 1351
rect 282 1348 334 1351
rect 338 1348 342 1351
rect 482 1348 502 1351
rect 506 1348 534 1351
rect 538 1348 782 1351
rect 858 1348 870 1351
rect 930 1348 1046 1351
rect 1050 1348 1070 1351
rect 1138 1348 1142 1351
rect 1146 1348 1161 1351
rect 1274 1348 1302 1351
rect 1342 1351 1345 1358
rect 1342 1348 1438 1351
rect 1594 1348 1654 1351
rect 1658 1348 1670 1351
rect 1714 1348 1782 1351
rect 110 1341 113 1348
rect 1158 1342 1161 1348
rect 1574 1342 1577 1348
rect 66 1338 113 1341
rect 314 1338 358 1341
rect 522 1338 534 1341
rect 562 1338 566 1341
rect 642 1338 726 1341
rect 954 1338 958 1341
rect 1026 1338 1030 1341
rect 1202 1338 1286 1341
rect 1474 1338 1534 1341
rect 1578 1338 1726 1341
rect 394 1328 414 1331
rect 434 1328 526 1331
rect 566 1331 569 1338
rect 566 1328 614 1331
rect 682 1328 710 1331
rect 826 1328 830 1331
rect 958 1331 961 1338
rect 958 1328 1014 1331
rect 1018 1328 1086 1331
rect 1194 1328 1238 1331
rect 1322 1328 1326 1331
rect 1330 1328 1350 1331
rect 1434 1328 1542 1331
rect 1666 1328 1670 1331
rect 1682 1328 1686 1331
rect 1698 1328 1782 1331
rect 1598 1322 1601 1328
rect 50 1318 62 1321
rect 66 1318 198 1321
rect 202 1318 374 1321
rect 498 1318 582 1321
rect 834 1318 878 1321
rect 898 1318 1406 1321
rect 1674 1318 1710 1321
rect 446 1312 449 1318
rect 734 1312 737 1318
rect 1478 1312 1481 1318
rect 66 1308 94 1311
rect 98 1308 230 1311
rect 818 1308 838 1311
rect 1154 1308 1294 1311
rect 1514 1308 1662 1311
rect 454 1302 457 1308
rect 888 1303 890 1307
rect 894 1303 897 1307
rect 902 1303 904 1307
rect 1038 1302 1041 1308
rect 514 1298 590 1301
rect 594 1298 638 1301
rect 674 1298 702 1301
rect 1082 1298 1102 1301
rect 1314 1298 1606 1301
rect 362 1288 430 1291
rect 434 1288 630 1291
rect 678 1288 758 1291
rect 1074 1288 1166 1291
rect 1170 1288 1270 1291
rect 1514 1288 1518 1291
rect 122 1278 222 1281
rect 354 1278 534 1281
rect 678 1281 681 1288
rect 606 1278 681 1281
rect 970 1278 1062 1281
rect 1238 1278 1310 1281
rect 1498 1278 1502 1281
rect 1634 1278 1646 1281
rect 1674 1278 1734 1281
rect 606 1272 609 1278
rect 686 1272 689 1278
rect 854 1272 857 1278
rect 298 1268 390 1271
rect 442 1268 454 1271
rect 530 1268 534 1271
rect 618 1268 638 1271
rect 642 1268 678 1271
rect 866 1268 958 1271
rect 1018 1268 1022 1271
rect 1158 1271 1161 1278
rect 1238 1272 1241 1278
rect 1342 1272 1345 1278
rect 1766 1272 1769 1278
rect 1158 1268 1206 1271
rect 1282 1268 1318 1271
rect 1350 1268 1358 1271
rect 1362 1268 1470 1271
rect 1642 1268 1686 1271
rect 26 1258 54 1261
rect 114 1258 161 1261
rect 394 1258 542 1261
rect 602 1258 606 1261
rect 654 1258 662 1261
rect 666 1258 726 1261
rect 794 1258 998 1261
rect 1034 1258 1062 1261
rect 1066 1258 1374 1261
rect 1686 1261 1689 1268
rect 1686 1258 1718 1261
rect 158 1252 161 1258
rect 1654 1252 1657 1258
rect 42 1248 102 1251
rect 218 1248 286 1251
rect 290 1248 438 1251
rect 442 1248 638 1251
rect 650 1248 718 1251
rect 746 1248 774 1251
rect 1002 1248 1006 1251
rect 1042 1248 1358 1251
rect 1362 1248 1614 1251
rect 1618 1248 1622 1251
rect 1662 1251 1665 1258
rect 1662 1248 1734 1251
rect 50 1238 158 1241
rect 258 1238 398 1241
rect 642 1238 646 1241
rect 650 1238 662 1241
rect 730 1238 1022 1241
rect 1026 1238 1142 1241
rect 1338 1238 1598 1241
rect 1706 1238 1798 1241
rect 402 1228 606 1231
rect 730 1228 990 1231
rect 994 1228 1150 1231
rect 1154 1228 1286 1231
rect 1298 1228 1334 1231
rect 378 1218 414 1221
rect 522 1218 766 1221
rect 1410 1218 1750 1221
rect 1798 1212 1801 1218
rect 970 1208 974 1211
rect 1626 1208 1670 1211
rect 368 1203 370 1207
rect 374 1203 377 1207
rect 382 1203 384 1207
rect 1384 1203 1386 1207
rect 1390 1203 1393 1207
rect 1398 1203 1400 1207
rect 74 1188 289 1191
rect 286 1181 289 1188
rect 286 1178 398 1181
rect 958 1181 961 1188
rect 958 1178 974 1181
rect 1618 1178 1670 1181
rect 1698 1178 1718 1181
rect 254 1172 257 1178
rect 26 1168 94 1171
rect 434 1168 502 1171
rect 722 1168 742 1171
rect 834 1168 942 1171
rect 954 1168 958 1171
rect 970 1168 990 1171
rect 1402 1168 1710 1171
rect 42 1158 78 1161
rect 82 1158 166 1161
rect 170 1158 318 1161
rect 322 1158 446 1161
rect 450 1158 478 1161
rect 642 1158 926 1161
rect 1126 1161 1129 1168
rect 1126 1158 1214 1161
rect 1330 1158 1574 1161
rect 1602 1158 1654 1161
rect 1694 1152 1697 1158
rect 26 1148 54 1151
rect 162 1148 366 1151
rect 474 1148 566 1151
rect 714 1148 726 1151
rect 754 1148 782 1151
rect 850 1148 854 1151
rect 914 1148 1046 1151
rect 1154 1148 1606 1151
rect 1150 1142 1153 1148
rect 186 1138 198 1141
rect 330 1138 350 1141
rect 426 1138 862 1141
rect 866 1138 982 1141
rect 986 1138 1070 1141
rect 1322 1138 1326 1141
rect 1362 1138 1462 1141
rect 1602 1138 1614 1141
rect 1626 1138 1630 1141
rect 1666 1138 1702 1141
rect 62 1131 65 1138
rect 62 1128 158 1131
rect 258 1128 342 1131
rect 354 1128 422 1131
rect 658 1128 694 1131
rect 762 1128 830 1131
rect 938 1128 966 1131
rect 1082 1128 1214 1131
rect 1362 1128 1438 1131
rect 1442 1128 1446 1131
rect 1450 1128 1526 1131
rect 1554 1128 1638 1131
rect 1650 1128 1734 1131
rect 234 1118 310 1121
rect 370 1118 470 1121
rect 818 1118 878 1121
rect 1018 1118 1094 1121
rect 1098 1118 1150 1121
rect 1378 1118 1470 1121
rect 1514 1118 1518 1121
rect 366 1111 369 1118
rect 314 1108 369 1111
rect 602 1108 630 1111
rect 994 1108 1070 1111
rect 1730 1108 1742 1111
rect 888 1103 890 1107
rect 894 1103 897 1107
rect 902 1103 904 1107
rect 546 1098 806 1101
rect 970 1098 990 1101
rect 1578 1098 1622 1101
rect 66 1088 126 1091
rect 130 1088 166 1091
rect 170 1088 246 1091
rect 250 1088 302 1091
rect 394 1088 462 1091
rect 1098 1088 1102 1091
rect 1626 1088 1686 1091
rect 210 1078 278 1081
rect 434 1078 550 1081
rect 562 1078 574 1081
rect 582 1078 974 1081
rect 986 1078 1318 1081
rect 1346 1078 1438 1081
rect 122 1068 134 1071
rect 138 1068 198 1071
rect 418 1068 422 1071
rect 466 1068 526 1071
rect 582 1071 585 1078
rect 1662 1072 1665 1078
rect 578 1068 585 1071
rect 778 1068 782 1071
rect 826 1068 838 1071
rect 866 1068 1070 1071
rect 1266 1068 1313 1071
rect 1434 1068 1462 1071
rect 1466 1068 1470 1071
rect 1482 1068 1494 1071
rect 1634 1068 1638 1071
rect 1690 1068 1702 1071
rect 1310 1062 1313 1068
rect 38 1058 126 1061
rect 226 1058 422 1061
rect 426 1058 614 1061
rect 642 1058 654 1061
rect 994 1058 998 1061
rect 1002 1058 1030 1061
rect 1130 1058 1158 1061
rect 1490 1058 1550 1061
rect 1554 1058 1601 1061
rect 1618 1058 1622 1061
rect 1646 1061 1649 1068
rect 1646 1058 1678 1061
rect 1682 1058 1694 1061
rect 1738 1058 1758 1061
rect 38 1052 41 1058
rect 1438 1052 1441 1058
rect 1598 1052 1601 1058
rect 330 1048 433 1051
rect 482 1048 510 1051
rect 562 1048 566 1051
rect 570 1048 606 1051
rect 642 1048 646 1051
rect 1658 1048 1670 1051
rect 1770 1048 1782 1051
rect 430 1042 433 1048
rect 410 1038 414 1041
rect 454 1038 510 1041
rect 650 1038 1006 1041
rect 1210 1038 1230 1041
rect 1794 1038 1798 1041
rect 278 1031 281 1038
rect 454 1031 457 1038
rect 278 1028 457 1031
rect 466 1028 486 1031
rect 498 1028 510 1031
rect 794 1028 1350 1031
rect 94 1021 97 1028
rect 94 1018 150 1021
rect 630 1021 633 1028
rect 330 1018 633 1021
rect 682 1018 830 1021
rect 858 1018 966 1021
rect 970 1018 1134 1021
rect 1290 1018 1294 1021
rect 1634 1018 1654 1021
rect 426 1008 478 1011
rect 618 1008 766 1011
rect 770 1008 982 1011
rect 986 1008 1334 1011
rect 1474 1008 1630 1011
rect 368 1003 370 1007
rect 374 1003 377 1007
rect 382 1003 384 1007
rect 1384 1003 1386 1007
rect 1390 1003 1393 1007
rect 1398 1003 1400 1007
rect 458 998 734 1001
rect 1538 998 1590 1001
rect 862 992 865 998
rect 162 988 422 991
rect 914 988 942 991
rect 946 988 998 991
rect 1338 988 1598 991
rect 1602 988 1646 991
rect 1142 982 1145 988
rect 138 978 182 981
rect 194 978 198 981
rect 202 978 406 981
rect 458 978 462 981
rect 506 978 878 981
rect 94 971 97 978
rect 94 968 358 971
rect 386 968 398 971
rect 402 968 486 971
rect 562 968 622 971
rect 650 968 766 971
rect 818 968 998 971
rect 1002 968 1046 971
rect 1486 962 1489 968
rect 154 958 166 961
rect 242 958 302 961
rect 338 958 366 961
rect 370 958 470 961
rect 474 958 478 961
rect 922 958 958 961
rect 962 958 966 961
rect 1330 958 1374 961
rect 1490 958 1534 961
rect 1606 961 1609 968
rect 1606 958 1710 961
rect 34 948 118 951
rect 130 948 142 951
rect 218 948 246 951
rect 298 948 422 951
rect 426 948 470 951
rect 474 948 598 951
rect 634 948 702 951
rect 734 951 737 958
rect 734 948 918 951
rect 1010 948 1062 951
rect 1074 948 1126 951
rect 1130 948 1134 951
rect 1226 948 1590 951
rect 1622 948 1638 951
rect 1582 942 1585 948
rect 1622 942 1625 948
rect 106 938 198 941
rect 202 938 254 941
rect 426 938 446 941
rect 458 938 462 941
rect 538 938 558 941
rect 738 938 806 941
rect 830 938 926 941
rect 970 938 1046 941
rect 1130 938 1150 941
rect 1154 938 1374 941
rect 830 932 833 938
rect 210 928 225 931
rect 250 928 318 931
rect 322 928 430 931
rect 458 928 558 931
rect 578 928 582 931
rect 962 928 982 931
rect 1178 928 1750 931
rect 222 922 225 928
rect 226 918 254 921
rect 410 918 422 921
rect 426 918 462 921
rect 554 918 598 921
rect 746 918 758 921
rect 762 918 998 921
rect 1162 918 1278 921
rect 1362 918 1430 921
rect 1474 918 1646 921
rect 1666 918 1734 921
rect 378 908 646 911
rect 1242 908 1294 911
rect 1410 908 1526 911
rect 1530 908 1774 911
rect 888 903 890 907
rect 894 903 897 907
rect 902 903 904 907
rect 122 898 214 901
rect 522 898 598 901
rect 706 898 750 901
rect 1002 898 1022 901
rect 1506 898 1510 901
rect 106 888 150 891
rect 258 888 286 891
rect 482 888 518 891
rect 538 888 590 891
rect 602 888 622 891
rect 626 888 830 891
rect 842 888 1150 891
rect 1482 888 1614 891
rect 1634 888 1638 891
rect 114 878 142 881
rect 178 878 206 881
rect 210 878 270 881
rect 274 878 433 881
rect 570 878 678 881
rect 698 878 934 881
rect 942 878 1022 881
rect 1450 878 1497 881
rect 1586 878 1638 881
rect 1670 881 1673 888
rect 1670 878 1710 881
rect 1730 878 1734 881
rect 1746 878 1798 881
rect 430 872 433 878
rect 202 868 222 871
rect 226 868 294 871
rect 434 868 438 871
rect 666 868 686 871
rect 942 871 945 878
rect 1494 872 1497 878
rect 850 868 945 871
rect 954 868 990 871
rect 1018 868 1062 871
rect 1594 868 1598 871
rect 1642 868 1782 871
rect 446 862 449 868
rect 34 858 102 861
rect 178 858 238 861
rect 258 858 262 861
rect 338 858 342 861
rect 354 858 438 861
rect 566 861 569 868
rect 774 862 777 868
rect 1166 862 1169 868
rect 482 858 569 861
rect 578 858 622 861
rect 626 858 657 861
rect 682 858 702 861
rect 834 858 958 861
rect 978 858 982 861
rect 994 858 1030 861
rect 1234 858 1254 861
rect 1666 858 1686 861
rect 1706 858 1710 861
rect 186 848 190 851
rect 282 848 406 851
rect 410 848 526 851
rect 642 848 646 851
rect 654 851 657 858
rect 654 848 950 851
rect 1162 848 1174 851
rect 1194 848 1230 851
rect 1378 848 1550 851
rect 1554 848 1622 851
rect 1626 848 1702 851
rect 1706 848 1718 851
rect 462 842 465 848
rect 218 838 238 841
rect 258 838 302 841
rect 354 838 390 841
rect 450 838 454 841
rect 650 838 694 841
rect 698 838 766 841
rect 810 838 870 841
rect 938 838 966 841
rect 970 838 1142 841
rect 1674 838 1750 841
rect 570 828 750 831
rect 278 822 281 828
rect 282 818 398 821
rect 402 818 430 821
rect 666 818 694 821
rect 722 818 742 821
rect 746 818 1006 821
rect 1322 818 1326 821
rect 762 808 1206 811
rect 1282 808 1334 811
rect 368 803 370 807
rect 374 803 377 807
rect 382 803 384 807
rect 394 798 534 801
rect 758 801 761 808
rect 1384 803 1386 807
rect 1390 803 1393 807
rect 1398 803 1400 807
rect 730 798 761 801
rect 1010 798 1326 801
rect 1330 798 1358 801
rect 266 788 745 791
rect 786 788 910 791
rect 1026 788 1110 791
rect 1114 788 1142 791
rect 1706 788 1710 791
rect 742 782 745 788
rect 202 778 222 781
rect 226 778 286 781
rect 394 778 438 781
rect 442 778 518 781
rect 634 778 734 781
rect 834 778 862 781
rect 866 778 974 781
rect 1026 778 1054 781
rect 1090 778 1142 781
rect 1146 778 1222 781
rect 1242 778 1390 781
rect 126 771 129 778
rect 126 768 238 771
rect 562 768 638 771
rect 738 768 870 771
rect 938 768 1006 771
rect 1010 768 1118 771
rect 1130 768 1134 771
rect 1186 768 1238 771
rect 1250 768 1286 771
rect 1314 768 1374 771
rect 194 758 209 761
rect 218 758 230 761
rect 454 758 494 761
rect 498 758 502 761
rect 554 758 614 761
rect 666 758 918 761
rect 922 758 1326 761
rect 34 748 158 751
rect 206 751 209 758
rect 454 752 457 758
rect 206 748 230 751
rect 306 748 374 751
rect 506 748 638 751
rect 698 748 750 751
rect 1002 748 1070 751
rect 1074 748 1142 751
rect 1146 748 1270 751
rect 1274 748 1286 751
rect 1298 748 1334 751
rect 1350 751 1353 758
rect 1430 752 1433 758
rect 1350 748 1422 751
rect 1578 748 1622 751
rect 1654 751 1657 758
rect 1626 748 1657 751
rect 1690 748 1750 751
rect 846 742 849 748
rect 98 738 142 741
rect 578 738 678 741
rect 826 738 830 741
rect 970 738 974 741
rect 1066 738 1438 741
rect 1442 738 1662 741
rect 1666 738 1742 741
rect 42 728 118 731
rect 154 728 206 731
rect 634 728 702 731
rect 1010 728 1022 731
rect 1026 728 1166 731
rect 1330 728 1406 731
rect 1450 728 1561 731
rect 1190 722 1193 728
rect 1558 722 1561 728
rect 66 718 158 721
rect 442 718 542 721
rect 546 718 598 721
rect 706 718 782 721
rect 818 718 854 721
rect 1106 718 1174 721
rect 1346 718 1470 721
rect 1638 718 1686 721
rect 1690 718 1758 721
rect 1638 712 1641 718
rect 578 708 774 711
rect 778 708 846 711
rect 954 708 998 711
rect 1042 708 1182 711
rect 1242 708 1382 711
rect 1386 708 1534 711
rect 888 703 890 707
rect 894 703 897 707
rect 902 703 904 707
rect 1550 702 1553 708
rect 90 698 102 701
rect 554 698 558 701
rect 650 698 726 701
rect 982 698 1102 701
rect 1106 698 1270 701
rect 982 692 985 698
rect 106 688 110 691
rect 186 688 286 691
rect 490 688 673 691
rect 802 688 862 691
rect 930 688 982 691
rect 1002 688 1014 691
rect 1082 688 1110 691
rect 1122 688 1414 691
rect 1546 688 1566 691
rect 1586 688 1638 691
rect 1646 688 1670 691
rect 670 682 673 688
rect 1646 682 1649 688
rect 258 678 262 681
rect 266 678 278 681
rect 290 678 486 681
rect 490 678 534 681
rect 538 678 566 681
rect 914 678 1017 681
rect 1014 672 1017 678
rect 1218 678 1358 681
rect 1442 678 1614 681
rect 1166 672 1169 678
rect 58 668 198 671
rect 226 668 262 671
rect 458 668 510 671
rect 546 668 550 671
rect 626 668 638 671
rect 730 668 854 671
rect 858 668 918 671
rect 986 668 998 671
rect 1034 668 1038 671
rect 1178 668 1214 671
rect 1242 668 1342 671
rect 1630 671 1633 678
rect 1418 668 1678 671
rect 82 658 142 661
rect 190 658 214 661
rect 242 658 326 661
rect 422 661 425 668
rect 678 662 681 668
rect 386 658 425 661
rect 434 658 494 661
rect 498 658 662 661
rect 746 658 814 661
rect 1070 661 1073 668
rect 874 658 1073 661
rect 1178 658 1182 661
rect 1234 658 1273 661
rect 1354 658 1358 661
rect 1410 658 1606 661
rect 1618 658 1646 661
rect 1682 658 1726 661
rect 190 652 193 658
rect 854 652 857 658
rect 862 652 865 658
rect 1270 652 1273 658
rect -26 651 -22 652
rect -26 648 6 651
rect 202 648 206 651
rect 602 648 830 651
rect 922 648 1054 651
rect 1058 648 1158 651
rect 1162 648 1198 651
rect 1434 648 1478 651
rect 1522 648 1526 651
rect 1554 648 1670 651
rect 1674 648 1686 651
rect 194 638 566 641
rect 610 638 726 641
rect 850 638 958 641
rect 962 638 1062 641
rect 1458 638 1462 641
rect 1602 638 1630 641
rect 434 628 438 631
rect 482 628 782 631
rect 1018 628 1038 631
rect 1378 628 1542 631
rect 642 618 718 621
rect 722 618 894 621
rect 1218 618 1422 621
rect 1434 618 1446 621
rect 1706 618 1710 621
rect 802 608 838 611
rect 858 608 1310 611
rect 1658 608 1694 611
rect 368 603 370 607
rect 374 603 377 607
rect 382 603 384 607
rect 1384 603 1386 607
rect 1390 603 1393 607
rect 1398 603 1400 607
rect 474 598 526 601
rect 778 598 838 601
rect 842 598 982 601
rect 1010 598 1014 601
rect 1018 598 1102 601
rect 1242 598 1366 601
rect 1426 598 1518 601
rect 1618 598 1638 601
rect 98 588 206 591
rect 210 588 238 591
rect 242 588 670 591
rect 674 588 1182 591
rect 1190 588 1574 591
rect 1578 588 1662 591
rect 1714 588 1766 591
rect 1190 582 1193 588
rect 1330 578 1422 581
rect 1482 578 1598 581
rect 50 568 222 571
rect 446 571 449 578
rect 1006 572 1009 578
rect 1790 572 1793 578
rect 446 568 462 571
rect 1154 568 1494 571
rect 1498 568 1574 571
rect 1578 568 1686 571
rect 74 558 134 561
rect 138 558 246 561
rect 278 561 281 568
rect 278 558 334 561
rect 498 558 502 561
rect 562 558 582 561
rect 586 558 622 561
rect 738 558 918 561
rect 1338 558 1361 561
rect 1394 558 1430 561
rect 1442 558 1638 561
rect 1642 558 1654 561
rect 1706 558 1798 561
rect 1190 552 1193 558
rect 26 548 54 551
rect 266 548 286 551
rect 306 548 406 551
rect 474 548 494 551
rect 522 548 542 551
rect 546 548 566 551
rect 786 548 942 551
rect 978 548 990 551
rect 222 542 225 548
rect 702 542 705 548
rect 1066 548 1118 551
rect 1138 548 1142 551
rect 1210 548 1302 551
rect 1358 551 1361 558
rect 1358 548 1382 551
rect 1410 548 1414 551
rect 1562 548 1582 551
rect 250 538 406 541
rect 410 538 678 541
rect 818 538 822 541
rect 970 538 998 541
rect 1242 538 1246 541
rect 1350 541 1353 548
rect 1766 542 1769 548
rect 1350 538 1422 541
rect 1426 538 1457 541
rect 1498 538 1558 541
rect 1618 538 1686 541
rect 30 532 33 538
rect 1454 532 1457 538
rect 66 528 166 531
rect 170 528 214 531
rect 218 528 318 531
rect 490 528 502 531
rect 514 528 614 531
rect 674 528 694 531
rect 738 528 758 531
rect 906 528 974 531
rect 562 518 622 521
rect 650 518 790 521
rect 794 518 806 521
rect 810 518 870 521
rect 882 518 1054 521
rect 1058 518 1102 521
rect 1282 518 1366 521
rect 1546 518 1750 521
rect 178 508 198 511
rect 202 508 446 511
rect 1034 508 1166 511
rect 1202 508 1438 511
rect 1538 508 1550 511
rect 1570 508 1614 511
rect 1738 508 1774 511
rect 888 503 890 507
rect 894 503 897 507
rect 902 503 904 507
rect 418 498 454 501
rect 458 498 534 501
rect 922 498 1078 501
rect 1186 498 1222 501
rect 94 491 97 498
rect 82 488 97 491
rect 354 488 438 491
rect 442 488 446 491
rect 602 488 678 491
rect 682 488 686 491
rect 914 488 974 491
rect 1086 488 1094 491
rect 1098 488 1214 491
rect 1218 488 1238 491
rect 1566 491 1569 498
rect 1562 488 1569 491
rect 1666 488 1678 491
rect 274 478 454 481
rect 618 478 718 481
rect 754 478 926 481
rect 986 478 1014 481
rect 1050 478 1086 481
rect 1090 478 1198 481
rect 1210 478 1366 481
rect 1466 478 1598 481
rect 166 471 169 478
rect 1662 472 1665 478
rect 1686 472 1689 478
rect 130 468 169 471
rect 530 468 537 471
rect 546 468 550 471
rect 658 468 686 471
rect 770 468 817 471
rect 842 468 934 471
rect 1130 468 1278 471
rect 1314 468 1334 471
rect 278 462 281 468
rect 170 458 230 461
rect 234 458 278 461
rect 382 461 385 468
rect 322 458 385 461
rect 534 461 537 468
rect 814 462 817 468
rect 534 458 598 461
rect 602 458 630 461
rect 874 458 974 461
rect 978 458 1030 461
rect 1130 458 1222 461
rect 1242 458 1270 461
rect 1342 461 1345 468
rect 1290 458 1345 461
rect 1598 461 1601 468
rect 1506 458 1694 461
rect 1722 458 1758 461
rect 90 448 190 451
rect 426 448 718 451
rect 818 448 822 451
rect 1170 448 1182 451
rect 1210 448 1246 451
rect 1322 448 1326 451
rect 1330 448 1478 451
rect 1546 448 1550 451
rect 1554 448 1670 451
rect 1698 448 1742 451
rect 1766 442 1769 448
rect 154 438 254 441
rect 258 438 358 441
rect 362 438 574 441
rect 882 438 894 441
rect 1370 438 1462 441
rect 1562 438 1582 441
rect 210 428 809 431
rect 818 428 1006 431
rect 1010 428 1046 431
rect 1050 428 1142 431
rect 202 418 286 421
rect 290 418 782 421
rect 806 421 809 428
rect 806 418 1486 421
rect 1490 418 1622 421
rect 1718 412 1721 418
rect 458 408 1326 411
rect 1610 408 1630 411
rect 1634 408 1646 411
rect 368 403 370 407
rect 374 403 377 407
rect 382 403 384 407
rect 1384 403 1386 407
rect 1390 403 1393 407
rect 1398 403 1400 407
rect 146 398 206 401
rect 450 398 534 401
rect 978 398 1014 401
rect 1522 398 1582 401
rect 1586 398 1670 401
rect 1722 398 1726 401
rect 654 388 702 391
rect 706 388 806 391
rect 946 388 990 391
rect 994 388 1030 391
rect 1410 388 1414 391
rect 654 382 657 388
rect 794 378 1062 381
rect 290 368 342 371
rect 346 368 462 371
rect 490 368 510 371
rect 554 368 558 371
rect 674 368 710 371
rect 714 368 750 371
rect 770 368 841 371
rect 890 368 918 371
rect 1050 368 1094 371
rect 1746 368 1782 371
rect 42 358 134 361
rect 282 358 286 361
rect 290 358 350 361
rect 542 361 545 368
rect 838 362 841 368
rect 410 358 545 361
rect 554 358 558 361
rect 650 358 654 361
rect 658 358 678 361
rect 706 358 726 361
rect 826 358 830 361
rect 910 358 974 361
rect 1010 358 1638 361
rect 50 348 102 351
rect 182 351 185 358
rect 910 352 913 358
rect 182 348 230 351
rect 234 348 582 351
rect 694 348 718 351
rect 778 348 822 351
rect 826 348 846 351
rect 1074 348 1153 351
rect 1162 348 1198 351
rect 1226 348 1230 351
rect 1618 348 1702 351
rect 1758 351 1761 358
rect 1754 348 1761 351
rect 226 338 302 341
rect 474 338 502 341
rect 506 338 529 341
rect 634 338 638 341
rect 686 341 689 348
rect 642 338 689 341
rect 694 342 697 348
rect 958 341 961 348
rect 882 338 961 341
rect 1066 338 1086 341
rect 1150 341 1153 348
rect 1150 338 1182 341
rect 1186 338 1206 341
rect 1274 338 1345 341
rect 1682 338 1702 341
rect 34 328 294 331
rect 298 328 318 331
rect 322 328 350 331
rect 422 331 425 338
rect 526 332 529 338
rect 1342 332 1345 338
rect 1710 332 1713 338
rect 370 328 494 331
rect 538 328 598 331
rect 602 328 686 331
rect 690 328 758 331
rect 802 328 814 331
rect 874 328 1038 331
rect 1078 328 1142 331
rect 1226 328 1230 331
rect 1078 322 1081 328
rect 194 318 438 321
rect 538 318 630 321
rect 642 318 694 321
rect 762 318 854 321
rect 858 318 990 321
rect 1234 318 1374 321
rect 1378 318 1390 321
rect 1394 318 1470 321
rect 1474 318 1534 321
rect 1594 318 1646 321
rect 1082 308 1166 311
rect 1170 308 1238 311
rect 1258 308 1430 311
rect 888 303 890 307
rect 894 303 897 307
rect 902 303 904 307
rect 98 298 174 301
rect 594 298 630 301
rect 658 298 742 301
rect 1698 298 1710 301
rect 66 288 182 291
rect 186 288 214 291
rect 218 288 286 291
rect 314 288 374 291
rect 554 288 646 291
rect 682 288 798 291
rect 826 288 830 291
rect 834 288 918 291
rect 930 288 1006 291
rect 1194 288 1302 291
rect 1442 288 1446 291
rect 1694 288 1798 291
rect 1694 282 1697 288
rect 162 278 174 281
rect 178 278 430 281
rect 602 278 622 281
rect 714 278 806 281
rect 1250 278 1262 281
rect 1698 278 1702 281
rect 130 268 150 271
rect 162 268 278 271
rect 434 268 454 271
rect 458 268 614 271
rect 706 268 750 271
rect 770 268 798 271
rect 890 268 958 271
rect 1218 268 1326 271
rect 1538 268 1734 271
rect 50 258 118 261
rect 210 258 406 261
rect 490 258 510 261
rect 514 258 550 261
rect 562 258 574 261
rect 578 258 598 261
rect 618 258 622 261
rect 626 258 630 261
rect 642 258 742 261
rect 746 258 974 261
rect 978 258 982 261
rect 1042 258 1110 261
rect 1146 258 1158 261
rect 1162 258 1270 261
rect 1274 258 1502 261
rect 1506 258 1582 261
rect 1586 258 1614 261
rect 1746 258 1790 261
rect 1302 252 1305 258
rect 34 248 38 251
rect 138 248 150 251
rect 154 248 230 251
rect 466 248 494 251
rect 498 248 678 251
rect 1146 248 1166 251
rect 1170 248 1238 251
rect 1466 248 1510 251
rect 1546 248 1734 251
rect 422 241 425 248
rect 1366 242 1369 248
rect 422 238 497 241
rect 610 238 750 241
rect 1690 238 1718 241
rect 494 232 497 238
rect 506 228 614 231
rect 850 228 1374 231
rect 1378 228 1414 231
rect 1418 228 1566 231
rect 1570 228 1694 231
rect 1722 228 1742 231
rect 346 218 374 221
rect 494 218 502 221
rect 506 218 510 221
rect 522 218 686 221
rect 1370 218 1454 221
rect 1698 218 1782 221
rect 970 208 998 211
rect 1002 208 1126 211
rect 1130 208 1182 211
rect 1186 208 1214 211
rect 368 203 370 207
rect 374 203 377 207
rect 382 203 384 207
rect 1384 203 1386 207
rect 1390 203 1393 207
rect 1398 203 1400 207
rect 754 198 878 201
rect 882 198 1118 201
rect 378 188 414 191
rect 802 188 806 191
rect 810 188 910 191
rect 978 188 982 191
rect 986 188 1070 191
rect 1622 191 1625 198
rect 1602 188 1625 191
rect 98 178 190 181
rect 1410 178 1526 181
rect 1530 178 1590 181
rect 1366 172 1369 178
rect 50 168 222 171
rect 282 168 670 171
rect 882 168 1006 171
rect 1410 168 1470 171
rect 1474 168 1486 171
rect 1550 168 1790 171
rect 18 158 54 161
rect 322 158 606 161
rect 690 158 790 161
rect 954 158 958 161
rect 1102 161 1105 168
rect 1042 158 1105 161
rect 1146 158 1158 161
rect 1178 158 1198 161
rect 1226 158 1286 161
rect 1550 161 1553 168
rect 1490 158 1553 161
rect 1666 158 1702 161
rect 1730 158 1758 161
rect 42 148 62 151
rect 82 148 110 151
rect 114 148 206 151
rect 226 148 390 151
rect 418 148 510 151
rect 514 148 654 151
rect 658 148 750 151
rect 862 151 865 158
rect 862 148 926 151
rect 954 148 1094 151
rect 1098 148 1174 151
rect 1210 148 1238 151
rect 1306 148 1382 151
rect 1486 151 1489 158
rect 1434 148 1489 151
rect 1558 151 1561 158
rect 1522 148 1561 151
rect 1650 148 1774 151
rect 1778 148 1782 151
rect 322 138 414 141
rect 530 138 534 141
rect 578 138 590 141
rect 594 138 718 141
rect 722 138 734 141
rect 738 138 1150 141
rect 1466 138 1478 141
rect 1482 138 1630 141
rect 130 128 166 131
rect 378 128 446 131
rect 494 131 497 138
rect 558 131 561 138
rect 1702 132 1705 138
rect 494 128 561 131
rect 570 128 598 131
rect 1178 128 1190 131
rect 1194 128 1198 131
rect 1410 128 1446 131
rect 1450 128 1494 131
rect 194 118 214 121
rect 1130 118 1238 121
rect 202 108 230 111
rect 1226 108 1230 111
rect 1642 108 1766 111
rect 888 103 890 107
rect 894 103 897 107
rect 902 103 904 107
rect 170 98 190 101
rect 970 98 1134 101
rect 1698 98 1718 101
rect 94 91 97 98
rect 1790 92 1793 98
rect 66 88 97 91
rect 282 88 334 91
rect 666 88 694 91
rect 1050 88 1118 91
rect 1122 88 1270 91
rect 1514 88 1606 91
rect 1610 88 1678 91
rect 162 78 222 81
rect 494 81 497 88
rect 418 78 497 81
rect 1202 78 1214 81
rect 1226 78 1230 81
rect 1298 78 1302 81
rect 1382 81 1385 88
rect 1362 78 1385 81
rect 1402 78 1406 81
rect 110 71 113 78
rect 58 68 113 71
rect 250 68 278 71
rect 374 71 377 78
rect 526 71 529 78
rect 298 68 529 71
rect 782 71 785 78
rect 1710 72 1713 78
rect 782 68 830 71
rect 906 68 1462 71
rect 1498 68 1534 71
rect 126 61 129 68
rect 90 58 129 61
rect 210 58 238 61
rect 242 58 262 61
rect 266 58 470 61
rect 474 58 502 61
rect 562 58 630 61
rect 718 61 721 68
rect 718 58 734 61
rect 778 58 862 61
rect 894 58 934 61
rect 1726 62 1729 68
rect 1026 59 1166 61
rect 1022 58 1166 59
rect 1226 58 1438 61
rect 1506 58 1510 61
rect 894 52 897 58
rect 202 48 894 51
rect 986 48 1470 51
rect 1082 38 1222 41
rect 570 8 574 11
rect 634 8 646 11
rect 778 8 790 11
rect 946 8 958 11
rect 368 3 370 7
rect 374 3 377 7
rect 382 3 384 7
rect 1384 3 1386 7
rect 1390 3 1393 7
rect 1398 3 1400 7
<< m4contact >>
rect 890 1703 894 1707
rect 898 1703 901 1707
rect 901 1703 902 1707
rect 518 1688 522 1692
rect 62 1658 66 1662
rect 406 1658 410 1662
rect 1038 1658 1042 1662
rect 1590 1658 1594 1662
rect 1646 1658 1650 1662
rect 1758 1658 1762 1662
rect 934 1648 938 1652
rect 446 1638 450 1642
rect 1014 1638 1018 1642
rect 1742 1638 1746 1642
rect 1782 1638 1786 1642
rect 1318 1628 1322 1632
rect 1694 1618 1698 1622
rect 1798 1618 1802 1622
rect 370 1603 374 1607
rect 378 1603 381 1607
rect 381 1603 382 1607
rect 1386 1603 1390 1607
rect 1394 1603 1397 1607
rect 1397 1603 1398 1607
rect 694 1598 698 1602
rect 1654 1598 1658 1602
rect 1790 1598 1794 1602
rect 878 1578 882 1582
rect 1798 1568 1802 1572
rect 598 1558 602 1562
rect 1678 1558 1682 1562
rect 1734 1558 1738 1562
rect 406 1548 410 1552
rect 766 1548 770 1552
rect 870 1548 874 1552
rect 1486 1548 1490 1552
rect 150 1538 154 1542
rect 1318 1538 1322 1542
rect 694 1518 698 1522
rect 1726 1518 1730 1522
rect 1006 1508 1010 1512
rect 890 1503 894 1507
rect 898 1503 901 1507
rect 901 1503 902 1507
rect 870 1498 874 1502
rect 1582 1478 1586 1482
rect 486 1468 490 1472
rect 622 1468 626 1472
rect 654 1468 658 1472
rect 854 1468 858 1472
rect 934 1468 938 1472
rect 1030 1468 1034 1472
rect 1558 1468 1562 1472
rect 1574 1468 1578 1472
rect 1686 1468 1690 1472
rect 774 1458 778 1462
rect 1006 1458 1010 1462
rect 1038 1458 1042 1462
rect 1342 1458 1346 1462
rect 1478 1458 1482 1462
rect 454 1448 458 1452
rect 462 1448 466 1452
rect 518 1418 522 1422
rect 686 1418 690 1422
rect 694 1408 698 1412
rect 1590 1408 1594 1412
rect 370 1403 374 1407
rect 378 1403 381 1407
rect 381 1403 382 1407
rect 1386 1403 1390 1407
rect 1394 1403 1397 1407
rect 1397 1403 1398 1407
rect 598 1388 602 1392
rect 998 1378 1002 1382
rect 646 1368 650 1372
rect 1038 1368 1042 1372
rect 1150 1368 1154 1372
rect 1750 1368 1754 1372
rect 230 1358 234 1362
rect 310 1358 314 1362
rect 574 1358 578 1362
rect 598 1358 602 1362
rect 342 1348 346 1352
rect 1134 1348 1138 1352
rect 1574 1348 1578 1352
rect 1590 1348 1594 1352
rect 1654 1348 1658 1352
rect 1710 1348 1714 1352
rect 534 1338 538 1342
rect 566 1338 570 1342
rect 638 1338 642 1342
rect 950 1338 954 1342
rect 1030 1338 1034 1342
rect 414 1328 418 1332
rect 830 1328 834 1332
rect 1326 1328 1330 1332
rect 1598 1328 1602 1332
rect 1662 1328 1666 1332
rect 1686 1328 1690 1332
rect 1694 1328 1698 1332
rect 62 1318 66 1322
rect 446 1318 450 1322
rect 830 1318 834 1322
rect 1478 1318 1482 1322
rect 1670 1318 1674 1322
rect 734 1308 738 1312
rect 1038 1308 1042 1312
rect 1662 1308 1666 1312
rect 890 1303 894 1307
rect 898 1303 901 1307
rect 901 1303 902 1307
rect 454 1298 458 1302
rect 686 1278 690 1282
rect 1342 1278 1346 1282
rect 1494 1278 1498 1282
rect 526 1268 530 1272
rect 854 1268 858 1272
rect 1014 1268 1018 1272
rect 1766 1268 1770 1272
rect 286 1248 290 1252
rect 638 1248 642 1252
rect 998 1248 1002 1252
rect 1614 1248 1618 1252
rect 1654 1248 1658 1252
rect 158 1238 162 1242
rect 398 1238 402 1242
rect 646 1238 650 1242
rect 726 1238 730 1242
rect 1702 1238 1706 1242
rect 1150 1228 1154 1232
rect 1798 1218 1802 1222
rect 974 1208 978 1212
rect 370 1203 374 1207
rect 378 1203 381 1207
rect 381 1203 382 1207
rect 1386 1203 1390 1207
rect 1394 1203 1397 1207
rect 1397 1203 1398 1207
rect 1718 1178 1722 1182
rect 254 1168 258 1172
rect 950 1168 954 1172
rect 478 1158 482 1162
rect 638 1158 642 1162
rect 1574 1158 1578 1162
rect 1694 1158 1698 1162
rect 726 1148 730 1152
rect 854 1148 858 1152
rect 1150 1148 1154 1152
rect 1606 1148 1610 1152
rect 1070 1138 1074 1142
rect 1318 1138 1322 1142
rect 1598 1138 1602 1142
rect 1622 1138 1626 1142
rect 1662 1138 1666 1142
rect 350 1128 354 1132
rect 310 1118 314 1122
rect 1518 1118 1522 1122
rect 1726 1108 1730 1112
rect 890 1103 894 1107
rect 898 1103 901 1107
rect 901 1103 902 1107
rect 966 1098 970 1102
rect 430 1078 434 1082
rect 1318 1078 1322 1082
rect 1662 1078 1666 1082
rect 422 1068 426 1072
rect 782 1068 786 1072
rect 838 1068 842 1072
rect 1470 1068 1474 1072
rect 222 1058 226 1062
rect 990 1058 994 1062
rect 1438 1058 1442 1062
rect 1614 1058 1618 1062
rect 1678 1058 1682 1062
rect 1734 1058 1738 1062
rect 558 1048 562 1052
rect 638 1048 642 1052
rect 1782 1048 1786 1052
rect 414 1038 418 1042
rect 1790 1038 1794 1042
rect 462 1028 466 1032
rect 854 1018 858 1022
rect 1134 1018 1138 1022
rect 1294 1018 1298 1022
rect 422 1008 426 1012
rect 766 1008 770 1012
rect 982 1008 986 1012
rect 1630 1008 1634 1012
rect 370 1003 374 1007
rect 378 1003 381 1007
rect 381 1003 382 1007
rect 1386 1003 1390 1007
rect 1394 1003 1397 1007
rect 1397 1003 1398 1007
rect 1534 998 1538 1002
rect 422 988 426 992
rect 862 988 866 992
rect 1646 988 1650 992
rect 190 978 194 982
rect 454 978 458 982
rect 1142 978 1146 982
rect 398 968 402 972
rect 558 968 562 972
rect 1486 968 1490 972
rect 334 958 338 962
rect 470 958 474 962
rect 734 958 738 962
rect 918 958 922 962
rect 598 948 602 952
rect 1006 948 1010 952
rect 1070 948 1074 952
rect 1134 948 1138 952
rect 1590 948 1594 952
rect 198 938 202 942
rect 454 938 458 942
rect 534 938 538 942
rect 1126 938 1130 942
rect 558 928 562 932
rect 574 928 578 932
rect 422 918 426 922
rect 462 918 466 922
rect 1470 918 1474 922
rect 1294 908 1298 912
rect 890 903 894 907
rect 898 903 901 907
rect 901 903 902 907
rect 1022 898 1026 902
rect 1502 898 1506 902
rect 598 888 602 892
rect 1150 888 1154 892
rect 1638 888 1642 892
rect 678 878 682 882
rect 934 878 938 882
rect 1734 878 1738 882
rect 1742 878 1746 882
rect 222 868 226 872
rect 430 868 434 872
rect 446 868 450 872
rect 774 868 778 872
rect 1166 868 1170 872
rect 1598 868 1602 872
rect 238 858 242 862
rect 254 858 258 862
rect 342 858 346 862
rect 438 858 442 862
rect 478 858 482 862
rect 982 858 986 862
rect 1662 858 1666 862
rect 1710 858 1714 862
rect 190 848 194 852
rect 638 848 642 852
rect 1550 848 1554 852
rect 454 838 458 842
rect 1750 838 1754 842
rect 750 828 754 832
rect 278 818 282 822
rect 370 803 374 807
rect 378 803 381 807
rect 381 803 382 807
rect 1386 803 1390 807
rect 1394 803 1397 807
rect 1397 803 1398 807
rect 1326 798 1330 802
rect 1702 788 1706 792
rect 286 778 290 782
rect 862 778 866 782
rect 1022 778 1026 782
rect 638 768 642 772
rect 870 768 874 772
rect 934 768 938 772
rect 1118 768 1122 772
rect 1126 768 1130 772
rect 230 758 234 762
rect 494 758 498 762
rect 1430 758 1434 762
rect 1142 748 1146 752
rect 1286 748 1290 752
rect 1334 748 1338 752
rect 1574 748 1578 752
rect 830 738 834 742
rect 846 738 850 742
rect 1438 738 1442 742
rect 1742 738 1746 742
rect 1166 728 1170 732
rect 1190 728 1194 732
rect 1406 728 1410 732
rect 702 718 706 722
rect 1174 718 1178 722
rect 1758 718 1762 722
rect 1534 708 1538 712
rect 1550 708 1554 712
rect 890 703 894 707
rect 898 703 901 707
rect 901 703 902 707
rect 550 698 554 702
rect 862 688 866 692
rect 1118 688 1122 692
rect 1566 688 1570 692
rect 1582 688 1586 692
rect 566 678 570 682
rect 1614 678 1618 682
rect 1646 678 1650 682
rect 542 668 546 672
rect 678 668 682 672
rect 726 668 730 672
rect 918 668 922 672
rect 998 668 1002 672
rect 1030 668 1034 672
rect 1166 668 1170 672
rect 854 658 858 662
rect 862 658 866 662
rect 870 658 874 662
rect 1174 658 1178 662
rect 1406 658 1410 662
rect 1614 658 1618 662
rect 206 648 210 652
rect 830 648 834 652
rect 1518 648 1522 652
rect 1686 648 1690 652
rect 726 638 730 642
rect 958 638 962 642
rect 1454 638 1458 642
rect 430 628 434 632
rect 782 628 786 632
rect 1014 628 1018 632
rect 638 618 642 622
rect 1422 618 1426 622
rect 1710 618 1714 622
rect 798 608 802 612
rect 1654 608 1658 612
rect 370 603 374 607
rect 378 603 381 607
rect 381 603 382 607
rect 1386 603 1390 607
rect 1394 603 1397 607
rect 1397 603 1398 607
rect 470 598 474 602
rect 1014 598 1018 602
rect 1422 598 1426 602
rect 1662 588 1666 592
rect 1766 588 1770 592
rect 1006 568 1010 572
rect 1790 568 1794 572
rect 494 558 498 562
rect 1190 558 1194 562
rect 1638 558 1642 562
rect 1798 558 1802 562
rect 702 548 706 552
rect 1134 548 1138 552
rect 1406 548 1410 552
rect 1582 548 1586 552
rect 1766 548 1770 552
rect 222 538 226 542
rect 406 538 410 542
rect 822 538 826 542
rect 1246 538 1250 542
rect 1494 538 1498 542
rect 30 528 34 532
rect 870 518 874 522
rect 1198 508 1202 512
rect 1734 508 1738 512
rect 890 503 894 507
rect 898 503 901 507
rect 901 503 902 507
rect 918 498 922 502
rect 446 488 450 492
rect 678 488 682 492
rect 1558 488 1562 492
rect 1678 488 1682 492
rect 750 478 754 482
rect 1198 478 1202 482
rect 1686 478 1690 482
rect 542 468 546 472
rect 1662 468 1666 472
rect 278 458 282 462
rect 870 458 874 462
rect 1126 458 1130 462
rect 1286 458 1290 462
rect 1718 458 1722 462
rect 422 448 426 452
rect 822 448 826 452
rect 1246 448 1250 452
rect 1318 448 1322 452
rect 1550 448 1554 452
rect 1670 448 1674 452
rect 1766 448 1770 452
rect 878 438 882 442
rect 1462 438 1466 442
rect 1142 428 1146 432
rect 198 418 202 422
rect 1606 408 1610 412
rect 1718 408 1722 412
rect 370 403 374 407
rect 378 403 381 407
rect 381 403 382 407
rect 1386 403 1390 407
rect 1394 403 1397 407
rect 1397 403 1398 407
rect 534 398 538 402
rect 974 398 978 402
rect 1726 398 1730 402
rect 702 388 706 392
rect 558 368 562 372
rect 766 368 770 372
rect 1742 368 1746 372
rect 1782 368 1786 372
rect 278 358 282 362
rect 558 358 562 362
rect 822 358 826 362
rect 230 348 234 352
rect 846 348 850 352
rect 1158 348 1162 352
rect 1230 348 1234 352
rect 1750 348 1754 352
rect 1182 338 1186 342
rect 1678 338 1682 342
rect 1710 338 1714 342
rect 30 328 34 332
rect 318 328 322 332
rect 350 328 354 332
rect 1230 328 1234 332
rect 630 318 634 322
rect 990 318 994 322
rect 1230 318 1234 322
rect 1166 308 1170 312
rect 890 303 894 307
rect 898 303 901 307
rect 901 303 902 307
rect 742 298 746 302
rect 1710 298 1714 302
rect 822 288 826 292
rect 1702 278 1706 282
rect 278 268 282 272
rect 574 258 578 262
rect 982 258 986 262
rect 30 248 34 252
rect 494 248 498 252
rect 1142 248 1146 252
rect 1366 248 1370 252
rect 1542 248 1546 252
rect 846 228 850 232
rect 1694 228 1698 232
rect 1718 228 1722 232
rect 370 203 374 207
rect 378 203 381 207
rect 381 203 382 207
rect 1386 203 1390 207
rect 1394 203 1397 207
rect 1397 203 1398 207
rect 878 198 882 202
rect 798 188 802 192
rect 974 188 978 192
rect 1366 178 1370 182
rect 278 168 282 172
rect 318 158 322 162
rect 950 158 954 162
rect 1158 158 1162 162
rect 1198 158 1202 162
rect 1286 158 1290 162
rect 1782 148 1786 152
rect 534 138 538 142
rect 1702 138 1706 142
rect 566 128 570 132
rect 1198 128 1202 132
rect 1406 128 1410 132
rect 1222 108 1226 112
rect 890 103 894 107
rect 898 103 901 107
rect 901 103 902 107
rect 1510 88 1514 92
rect 1790 88 1794 92
rect 1222 78 1226 82
rect 1302 78 1306 82
rect 1398 78 1402 82
rect 1710 68 1714 72
rect 1510 58 1514 62
rect 1726 58 1730 62
rect 982 48 986 52
rect 1222 38 1226 42
rect 574 8 578 12
rect 370 3 374 7
rect 378 3 381 7
rect 381 3 382 7
rect 1386 3 1390 7
rect 1394 3 1397 7
rect 1397 3 1398 7
<< metal4 >>
rect 888 1703 890 1707
rect 894 1703 897 1707
rect 902 1703 904 1707
rect 62 1322 65 1658
rect 368 1603 370 1607
rect 374 1603 377 1607
rect 382 1603 384 1607
rect 406 1552 409 1658
rect 154 1538 161 1541
rect 158 1242 161 1538
rect 368 1403 370 1407
rect 374 1403 377 1407
rect 382 1403 384 1407
rect 222 1358 230 1361
rect 222 1062 225 1358
rect 190 852 193 978
rect 198 651 201 938
rect 198 648 206 651
rect 30 332 33 528
rect 198 422 201 648
rect 222 542 225 868
rect 254 862 257 1168
rect 242 858 246 861
rect 230 352 233 758
rect 278 462 281 818
rect 286 782 289 1248
rect 310 1122 313 1358
rect 334 1348 342 1351
rect 334 962 337 1348
rect 342 1342 345 1348
rect 418 1328 422 1331
rect 446 1322 449 1638
rect 490 1468 494 1471
rect 454 1452 457 1468
rect 368 1203 370 1207
rect 374 1203 377 1207
rect 382 1203 384 1207
rect 338 858 342 861
rect 286 361 289 778
rect 282 358 289 361
rect 30 252 33 328
rect 278 272 281 358
rect 350 332 353 1128
rect 368 1003 370 1007
rect 374 1003 377 1007
rect 382 1003 384 1007
rect 398 972 401 1238
rect 406 1038 414 1041
rect 368 803 370 807
rect 374 803 377 807
rect 382 803 384 807
rect 368 603 370 607
rect 374 603 377 607
rect 382 603 384 607
rect 406 542 409 1038
rect 422 1012 425 1068
rect 422 992 425 1008
rect 422 452 425 918
rect 430 872 433 1078
rect 454 982 457 1298
rect 462 1032 465 1448
rect 518 1422 521 1688
rect 598 1392 601 1558
rect 694 1522 697 1598
rect 626 1468 633 1471
rect 658 1468 662 1471
rect 594 1358 598 1361
rect 562 1338 566 1341
rect 534 1271 537 1338
rect 530 1268 537 1271
rect 430 632 433 868
rect 438 862 441 868
rect 446 492 449 868
rect 454 842 457 938
rect 462 922 465 1028
rect 470 602 473 958
rect 478 862 481 1158
rect 562 1048 569 1051
rect 494 562 497 758
rect 368 403 370 407
rect 374 403 377 407
rect 382 403 384 407
rect 278 172 281 268
rect 318 162 321 328
rect 494 252 497 558
rect 534 402 537 938
rect 558 932 561 968
rect 542 472 545 668
rect 550 361 553 698
rect 566 682 569 1048
rect 574 932 577 1358
rect 598 892 601 948
rect 562 368 566 371
rect 550 358 558 361
rect 630 322 633 1468
rect 638 1252 641 1338
rect 646 1242 649 1368
rect 686 1282 689 1418
rect 694 1412 697 1518
rect 638 1052 641 1158
rect 726 1152 729 1238
rect 638 852 641 1048
rect 734 962 737 1308
rect 766 1012 769 1548
rect 870 1502 873 1548
rect 682 878 686 881
rect 774 872 777 1458
rect 826 1328 830 1331
rect 638 772 641 848
rect 638 622 641 768
rect 678 492 681 668
rect 702 552 705 718
rect 726 642 729 668
rect 702 392 705 548
rect 750 482 753 828
rect 782 632 785 1068
rect 830 742 833 1318
rect 854 1272 857 1468
rect 842 1068 846 1071
rect 854 1022 857 1148
rect 834 648 838 651
rect 762 368 766 371
rect 742 302 745 328
rect 368 203 370 207
rect 374 203 377 207
rect 382 203 384 207
rect 530 138 534 141
rect 566 132 569 138
rect 574 12 577 258
rect 798 192 801 608
rect 822 452 825 538
rect 822 292 825 358
rect 846 352 849 738
rect 854 662 857 1018
rect 862 782 865 988
rect 862 662 865 688
rect 870 662 873 768
rect 870 462 873 518
rect 878 442 881 1578
rect 888 1503 890 1507
rect 894 1503 897 1507
rect 902 1503 904 1507
rect 934 1472 937 1648
rect 1006 1638 1014 1641
rect 1006 1512 1009 1638
rect 1002 1458 1006 1461
rect 888 1303 890 1307
rect 894 1303 897 1307
rect 902 1303 904 1307
rect 950 1172 953 1338
rect 998 1252 1001 1378
rect 1030 1342 1033 1468
rect 1038 1462 1041 1658
rect 1318 1542 1321 1628
rect 1384 1603 1386 1607
rect 1390 1603 1393 1607
rect 1398 1603 1400 1607
rect 1038 1312 1041 1368
rect 966 1208 974 1211
rect 888 1103 890 1107
rect 894 1103 897 1107
rect 902 1103 904 1107
rect 966 1102 969 1208
rect 888 903 890 907
rect 894 903 897 907
rect 902 903 904 907
rect 888 703 890 707
rect 894 703 897 707
rect 902 703 904 707
rect 918 672 921 958
rect 934 772 937 878
rect 982 862 985 1008
rect 888 503 890 507
rect 894 503 897 507
rect 902 503 904 507
rect 918 502 921 668
rect 846 232 849 348
rect 878 202 881 438
rect 888 303 890 307
rect 894 303 897 307
rect 902 303 904 307
rect 958 161 961 638
rect 974 192 977 398
rect 982 262 985 858
rect 990 322 993 1058
rect 998 672 1001 678
rect 1006 601 1009 948
rect 1014 632 1017 1268
rect 1070 952 1073 1138
rect 1134 1022 1137 1348
rect 1150 1232 1153 1368
rect 1022 782 1025 898
rect 1126 772 1129 938
rect 1118 692 1121 768
rect 1026 668 1030 671
rect 1006 598 1014 601
rect 1006 572 1009 578
rect 1126 462 1129 768
rect 1134 552 1137 948
rect 1142 752 1145 978
rect 1150 892 1153 1148
rect 1318 1142 1321 1538
rect 1318 1082 1321 1138
rect 1294 912 1297 1018
rect 1162 868 1166 871
rect 1166 672 1169 728
rect 954 158 961 161
rect 888 103 890 107
rect 894 103 897 107
rect 902 103 904 107
rect 982 52 985 258
rect 1142 252 1145 428
rect 1158 162 1161 348
rect 1166 312 1169 668
rect 1174 662 1177 718
rect 1178 658 1185 661
rect 1182 342 1185 658
rect 1190 562 1193 728
rect 1198 482 1201 508
rect 1246 452 1249 538
rect 1286 462 1289 748
rect 1222 348 1230 351
rect 1198 132 1201 158
rect 1222 112 1225 348
rect 1230 322 1233 328
rect 1286 162 1289 458
rect 1318 452 1321 1078
rect 1326 802 1329 1328
rect 1342 1282 1345 1458
rect 1384 1403 1386 1407
rect 1390 1403 1393 1407
rect 1398 1403 1400 1407
rect 1478 1322 1481 1458
rect 1384 1203 1386 1207
rect 1390 1203 1393 1207
rect 1398 1203 1400 1207
rect 1384 1003 1386 1007
rect 1390 1003 1393 1007
rect 1398 1003 1400 1007
rect 1384 803 1386 807
rect 1390 803 1393 807
rect 1398 803 1400 807
rect 1430 752 1433 758
rect 1338 748 1342 751
rect 1438 742 1441 1058
rect 1470 922 1473 1068
rect 1486 972 1489 1548
rect 1570 1468 1574 1471
rect 1406 662 1409 728
rect 1384 603 1386 607
rect 1390 603 1393 607
rect 1398 603 1400 607
rect 1406 552 1409 658
rect 1458 638 1465 641
rect 1422 602 1425 618
rect 1384 403 1386 407
rect 1390 403 1393 407
rect 1398 403 1400 407
rect 1366 182 1369 248
rect 1384 203 1386 207
rect 1390 203 1393 207
rect 1398 203 1400 207
rect 1406 132 1409 548
rect 1462 442 1465 638
rect 1494 542 1497 1278
rect 1510 1118 1518 1121
rect 1298 78 1302 81
rect 1394 78 1398 81
rect 1222 42 1225 78
rect 1502 61 1505 898
rect 1510 92 1513 1118
rect 1534 712 1537 998
rect 1550 712 1553 848
rect 1522 648 1526 651
rect 1558 492 1561 1468
rect 1574 1162 1577 1348
rect 1574 752 1577 1158
rect 1582 692 1585 1478
rect 1590 1412 1593 1658
rect 1590 952 1593 1348
rect 1598 1142 1601 1328
rect 1598 872 1601 878
rect 1570 688 1574 691
rect 1582 552 1585 688
rect 1542 448 1550 451
rect 1542 252 1545 448
rect 1606 412 1609 1148
rect 1614 1062 1617 1248
rect 1626 1138 1633 1141
rect 1630 1012 1633 1138
rect 1646 992 1649 1658
rect 1654 1352 1657 1598
rect 1662 1312 1665 1328
rect 1614 662 1617 678
rect 1638 562 1641 888
rect 1646 682 1649 688
rect 1654 612 1657 1248
rect 1662 1142 1665 1308
rect 1662 1072 1665 1078
rect 1662 592 1665 858
rect 1662 472 1665 588
rect 1670 452 1673 1318
rect 1678 1062 1681 1558
rect 1686 1332 1689 1468
rect 1694 1332 1697 1618
rect 1678 342 1681 488
rect 1686 482 1689 648
rect 1694 232 1697 1158
rect 1702 792 1705 1238
rect 1710 862 1713 1348
rect 1710 342 1713 618
rect 1718 462 1721 1178
rect 1726 1132 1729 1518
rect 1702 142 1705 278
rect 1710 72 1713 298
rect 1718 232 1721 408
rect 1726 402 1729 1108
rect 1734 1062 1737 1558
rect 1742 882 1745 1638
rect 1734 512 1737 878
rect 1750 842 1753 1368
rect 1742 372 1745 738
rect 1750 352 1753 838
rect 1758 722 1761 1658
rect 1766 592 1769 1268
rect 1782 1052 1785 1638
rect 1790 1042 1793 1598
rect 1798 1572 1801 1618
rect 1766 452 1769 548
rect 1782 152 1785 368
rect 1790 92 1793 568
rect 1798 562 1801 1218
rect 1502 58 1510 61
rect 1722 58 1726 61
rect 368 3 370 7
rect 374 3 377 7
rect 382 3 384 7
rect 1384 3 1386 7
rect 1390 3 1393 7
rect 1398 3 1400 7
<< m5contact >>
rect 890 1703 894 1707
rect 897 1703 898 1707
rect 898 1703 901 1707
rect 370 1603 374 1607
rect 377 1603 378 1607
rect 378 1603 381 1607
rect 370 1403 374 1407
rect 377 1403 378 1407
rect 378 1403 381 1407
rect 310 1358 314 1362
rect 246 858 250 862
rect 342 1338 346 1342
rect 422 1328 426 1332
rect 454 1468 458 1472
rect 494 1468 498 1472
rect 370 1203 374 1207
rect 377 1203 378 1207
rect 378 1203 381 1207
rect 334 858 338 862
rect 370 1003 374 1007
rect 377 1003 378 1007
rect 378 1003 381 1007
rect 370 803 374 807
rect 377 803 378 807
rect 378 803 381 807
rect 370 603 374 607
rect 377 603 378 607
rect 378 603 381 607
rect 662 1468 666 1472
rect 590 1358 594 1362
rect 558 1338 562 1342
rect 438 868 442 872
rect 370 403 374 407
rect 377 403 378 407
rect 378 403 381 407
rect 566 368 570 372
rect 686 878 690 882
rect 822 1328 826 1332
rect 846 1068 850 1072
rect 838 648 842 652
rect 758 368 762 372
rect 742 328 746 332
rect 370 203 374 207
rect 377 203 378 207
rect 378 203 381 207
rect 526 138 530 142
rect 566 138 570 142
rect 890 1503 894 1507
rect 897 1503 898 1507
rect 898 1503 901 1507
rect 998 1458 1002 1462
rect 890 1303 894 1307
rect 897 1303 898 1307
rect 898 1303 901 1307
rect 1386 1603 1390 1607
rect 1393 1603 1394 1607
rect 1394 1603 1397 1607
rect 890 1103 894 1107
rect 897 1103 898 1107
rect 898 1103 901 1107
rect 890 903 894 907
rect 897 903 898 907
rect 898 903 901 907
rect 890 703 894 707
rect 897 703 898 707
rect 898 703 901 707
rect 890 503 894 507
rect 897 503 898 507
rect 898 503 901 507
rect 890 303 894 307
rect 897 303 898 307
rect 898 303 901 307
rect 998 678 1002 682
rect 1022 668 1026 672
rect 1006 578 1010 582
rect 1158 868 1162 872
rect 890 103 894 107
rect 897 103 898 107
rect 898 103 901 107
rect 1230 318 1234 322
rect 1386 1403 1390 1407
rect 1393 1403 1394 1407
rect 1394 1403 1397 1407
rect 1386 1203 1390 1207
rect 1393 1203 1394 1207
rect 1394 1203 1397 1207
rect 1386 1003 1390 1007
rect 1393 1003 1394 1007
rect 1394 1003 1397 1007
rect 1386 803 1390 807
rect 1393 803 1394 807
rect 1394 803 1397 807
rect 1342 748 1346 752
rect 1430 748 1434 752
rect 1566 1468 1570 1472
rect 1386 603 1390 607
rect 1393 603 1394 607
rect 1394 603 1397 607
rect 1386 403 1390 407
rect 1393 403 1394 407
rect 1394 403 1397 407
rect 1386 203 1390 207
rect 1393 203 1394 207
rect 1394 203 1397 207
rect 1294 78 1298 82
rect 1390 78 1394 82
rect 1526 648 1530 652
rect 1598 878 1602 882
rect 1574 688 1578 692
rect 1646 688 1650 692
rect 1662 1068 1666 1072
rect 1726 1128 1730 1132
rect 1718 58 1722 62
rect 370 3 374 7
rect 377 3 378 7
rect 378 3 381 7
rect 1386 3 1390 7
rect 1393 3 1394 7
rect 1394 3 1397 7
<< metal5 >>
rect 894 1703 897 1707
rect 893 1702 898 1703
rect 903 1702 904 1707
rect 374 1603 377 1607
rect 373 1602 378 1603
rect 383 1602 384 1607
rect 1390 1603 1393 1607
rect 1389 1602 1394 1603
rect 1399 1602 1400 1607
rect 894 1503 897 1507
rect 893 1502 898 1503
rect 903 1502 904 1507
rect 458 1468 494 1471
rect 666 1468 1566 1471
rect 1002 1458 1005 1461
rect 374 1403 377 1407
rect 373 1402 378 1403
rect 383 1402 384 1407
rect 1390 1403 1393 1407
rect 1389 1402 1394 1403
rect 1399 1402 1400 1407
rect 314 1358 590 1361
rect 346 1338 558 1341
rect 426 1328 822 1331
rect 894 1303 897 1307
rect 893 1302 898 1303
rect 903 1302 904 1307
rect 374 1203 377 1207
rect 373 1202 378 1203
rect 383 1202 384 1207
rect 1390 1203 1393 1207
rect 1389 1202 1394 1203
rect 1399 1202 1400 1207
rect 1726 1122 1729 1128
rect 894 1103 897 1107
rect 893 1102 898 1103
rect 903 1102 904 1107
rect 850 1068 1662 1071
rect 374 1003 377 1007
rect 373 1002 378 1003
rect 383 1002 384 1007
rect 1390 1003 1393 1007
rect 1389 1002 1394 1003
rect 1399 1002 1400 1007
rect 894 903 897 907
rect 893 902 898 903
rect 903 902 904 907
rect 690 878 1598 881
rect 442 868 1158 871
rect 250 858 334 861
rect 374 803 377 807
rect 373 802 378 803
rect 383 802 384 807
rect 1390 803 1393 807
rect 1389 802 1394 803
rect 1399 802 1400 807
rect 1346 748 1430 751
rect 894 703 897 707
rect 893 702 898 703
rect 903 702 904 707
rect 1578 688 1646 691
rect 998 671 1001 678
rect 998 668 1022 671
rect 842 648 1526 651
rect 374 603 377 607
rect 373 602 378 603
rect 383 602 384 607
rect 1390 603 1393 607
rect 1389 602 1394 603
rect 1399 602 1400 607
rect 1006 582 1009 587
rect 894 503 897 507
rect 893 502 898 503
rect 903 502 904 507
rect 374 403 377 407
rect 373 402 378 403
rect 383 402 384 407
rect 1390 403 1393 407
rect 1389 402 1394 403
rect 1399 402 1400 407
rect 570 368 758 371
rect 746 328 1233 331
rect 1230 322 1233 328
rect 894 303 897 307
rect 893 302 898 303
rect 903 302 904 307
rect 374 203 377 207
rect 373 202 378 203
rect 383 202 384 207
rect 1390 203 1393 207
rect 1389 202 1394 203
rect 1399 202 1400 207
rect 530 138 566 141
rect 894 103 897 107
rect 893 102 898 103
rect 903 102 904 107
rect 1298 78 1390 81
rect 1722 58 1725 61
rect 374 3 377 7
rect 373 2 378 3
rect 383 2 384 7
rect 1390 3 1393 7
rect 1389 2 1394 3
rect 1399 2 1400 7
<< m6contact >>
rect 888 1703 890 1707
rect 890 1703 893 1707
rect 898 1703 901 1707
rect 901 1703 903 1707
rect 888 1702 893 1703
rect 898 1702 903 1703
rect 368 1603 370 1607
rect 370 1603 373 1607
rect 378 1603 381 1607
rect 381 1603 383 1607
rect 368 1602 373 1603
rect 378 1602 383 1603
rect 1384 1603 1386 1607
rect 1386 1603 1389 1607
rect 1394 1603 1397 1607
rect 1397 1603 1399 1607
rect 1384 1602 1389 1603
rect 1394 1602 1399 1603
rect 888 1503 890 1507
rect 890 1503 893 1507
rect 898 1503 901 1507
rect 901 1503 903 1507
rect 888 1502 893 1503
rect 898 1502 903 1503
rect 1005 1457 1010 1462
rect 368 1403 370 1407
rect 370 1403 373 1407
rect 378 1403 381 1407
rect 381 1403 383 1407
rect 368 1402 373 1403
rect 378 1402 383 1403
rect 1384 1403 1386 1407
rect 1386 1403 1389 1407
rect 1394 1403 1397 1407
rect 1397 1403 1399 1407
rect 1384 1402 1389 1403
rect 1394 1402 1399 1403
rect 888 1303 890 1307
rect 890 1303 893 1307
rect 898 1303 901 1307
rect 901 1303 903 1307
rect 888 1302 893 1303
rect 898 1302 903 1303
rect 368 1203 370 1207
rect 370 1203 373 1207
rect 378 1203 381 1207
rect 381 1203 383 1207
rect 368 1202 373 1203
rect 378 1202 383 1203
rect 1384 1203 1386 1207
rect 1386 1203 1389 1207
rect 1394 1203 1397 1207
rect 1397 1203 1399 1207
rect 1384 1202 1389 1203
rect 1394 1202 1399 1203
rect 1725 1117 1730 1122
rect 888 1103 890 1107
rect 890 1103 893 1107
rect 898 1103 901 1107
rect 901 1103 903 1107
rect 888 1102 893 1103
rect 898 1102 903 1103
rect 368 1003 370 1007
rect 370 1003 373 1007
rect 378 1003 381 1007
rect 381 1003 383 1007
rect 368 1002 373 1003
rect 378 1002 383 1003
rect 1384 1003 1386 1007
rect 1386 1003 1389 1007
rect 1394 1003 1397 1007
rect 1397 1003 1399 1007
rect 1384 1002 1389 1003
rect 1394 1002 1399 1003
rect 888 903 890 907
rect 890 903 893 907
rect 898 903 901 907
rect 901 903 903 907
rect 888 902 893 903
rect 898 902 903 903
rect 368 803 370 807
rect 370 803 373 807
rect 378 803 381 807
rect 381 803 383 807
rect 368 802 373 803
rect 378 802 383 803
rect 1384 803 1386 807
rect 1386 803 1389 807
rect 1394 803 1397 807
rect 1397 803 1399 807
rect 1384 802 1389 803
rect 1394 802 1399 803
rect 888 703 890 707
rect 890 703 893 707
rect 898 703 901 707
rect 901 703 903 707
rect 888 702 893 703
rect 898 702 903 703
rect 368 603 370 607
rect 370 603 373 607
rect 378 603 381 607
rect 381 603 383 607
rect 368 602 373 603
rect 378 602 383 603
rect 1384 603 1386 607
rect 1386 603 1389 607
rect 1394 603 1397 607
rect 1397 603 1399 607
rect 1384 602 1389 603
rect 1394 602 1399 603
rect 1005 587 1010 592
rect 888 503 890 507
rect 890 503 893 507
rect 898 503 901 507
rect 901 503 903 507
rect 888 502 893 503
rect 898 502 903 503
rect 368 403 370 407
rect 370 403 373 407
rect 378 403 381 407
rect 381 403 383 407
rect 368 402 373 403
rect 378 402 383 403
rect 1384 403 1386 407
rect 1386 403 1389 407
rect 1394 403 1397 407
rect 1397 403 1399 407
rect 1384 402 1389 403
rect 1394 402 1399 403
rect 888 303 890 307
rect 890 303 893 307
rect 898 303 901 307
rect 901 303 903 307
rect 888 302 893 303
rect 898 302 903 303
rect 368 203 370 207
rect 370 203 373 207
rect 378 203 381 207
rect 381 203 383 207
rect 368 202 373 203
rect 378 202 383 203
rect 1384 203 1386 207
rect 1386 203 1389 207
rect 1394 203 1397 207
rect 1397 203 1399 207
rect 1384 202 1389 203
rect 1394 202 1399 203
rect 888 103 890 107
rect 890 103 893 107
rect 898 103 901 107
rect 901 103 903 107
rect 888 102 893 103
rect 898 102 903 103
rect 1725 57 1730 62
rect 368 3 370 7
rect 370 3 373 7
rect 378 3 381 7
rect 381 3 383 7
rect 368 2 373 3
rect 378 2 383 3
rect 1384 3 1386 7
rect 1386 3 1389 7
rect 1394 3 1397 7
rect 1397 3 1399 7
rect 1384 2 1389 3
rect 1394 2 1399 3
<< metal6 >>
rect 368 1607 384 1730
rect 373 1602 378 1607
rect 383 1602 384 1607
rect 368 1407 384 1602
rect 373 1402 378 1407
rect 383 1402 384 1407
rect 368 1207 384 1402
rect 373 1202 378 1207
rect 383 1202 384 1207
rect 368 1007 384 1202
rect 373 1002 378 1007
rect 383 1002 384 1007
rect 368 807 384 1002
rect 373 802 378 807
rect 383 802 384 807
rect 368 607 384 802
rect 373 602 378 607
rect 383 602 384 607
rect 368 407 384 602
rect 373 402 378 407
rect 383 402 384 407
rect 368 207 384 402
rect 373 202 378 207
rect 383 202 384 207
rect 368 7 384 202
rect 373 2 378 7
rect 383 2 384 7
rect 368 -30 384 2
rect 888 1707 904 1730
rect 893 1702 898 1707
rect 903 1702 904 1707
rect 888 1507 904 1702
rect 893 1502 898 1507
rect 903 1502 904 1507
rect 888 1307 904 1502
rect 1384 1607 1400 1730
rect 1389 1602 1394 1607
rect 1399 1602 1400 1607
rect 893 1302 898 1307
rect 903 1302 904 1307
rect 888 1107 904 1302
rect 893 1102 898 1107
rect 903 1102 904 1107
rect 888 907 904 1102
rect 893 902 898 907
rect 903 902 904 907
rect 888 707 904 902
rect 893 702 898 707
rect 903 702 904 707
rect 888 507 904 702
rect 1005 592 1010 1457
rect 1384 1407 1400 1602
rect 1389 1402 1394 1407
rect 1399 1402 1400 1407
rect 1384 1207 1400 1402
rect 1389 1202 1394 1207
rect 1399 1202 1400 1207
rect 1384 1007 1400 1202
rect 1389 1002 1394 1007
rect 1399 1002 1400 1007
rect 1384 807 1400 1002
rect 1389 802 1394 807
rect 1399 802 1400 807
rect 1384 607 1400 802
rect 1389 602 1394 607
rect 1399 602 1400 607
rect 893 502 898 507
rect 903 502 904 507
rect 888 307 904 502
rect 893 302 898 307
rect 903 302 904 307
rect 888 107 904 302
rect 893 102 898 107
rect 903 102 904 107
rect 888 -30 904 102
rect 1384 407 1400 602
rect 1389 402 1394 407
rect 1399 402 1400 407
rect 1384 207 1400 402
rect 1389 202 1394 207
rect 1399 202 1400 207
rect 1384 7 1400 202
rect 1725 62 1730 1117
rect 1389 2 1394 7
rect 1399 2 1400 7
rect 1384 -30 1400 2
use DFFPOSX1  DFFPOSX1_7
timestamp 1751994658
transform 1 0 4 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1751994658
transform 1 0 100 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_16
timestamp 1751994658
transform -1 0 52 0 1 105
box -2 -3 50 103
use INVX1  INVX1_17
timestamp 1751994658
transform -1 0 68 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_15
timestamp 1751994658
transform 1 0 68 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_26
timestamp 1751994658
transform -1 0 124 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1751994658
transform -1 0 220 0 1 105
box -2 -3 98 103
use AOI21X1  AOI21X1_16
timestamp 1751994658
transform 1 0 196 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1751994658
transform 1 0 228 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1751994658
transform 1 0 252 0 -1 105
box -2 -3 98 103
use FILL  FILL_0_0_0
timestamp 1751994658
transform 1 0 348 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1751994658
transform 1 0 356 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1751994658
transform 1 0 364 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_17
timestamp 1751994658
transform 1 0 220 0 1 105
box -2 -3 50 103
use INVX1  INVX1_18
timestamp 1751994658
transform -1 0 284 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1751994658
transform 1 0 284 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_23
timestamp 1751994658
transform 1 0 460 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1751994658
transform -1 0 516 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1751994658
transform 1 0 516 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_0_0
timestamp 1751994658
transform 1 0 380 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1751994658
transform 1 0 388 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_13
timestamp 1751994658
transform 1 0 396 0 1 105
box -2 -3 50 103
use INVX1  INVX1_14
timestamp 1751994658
transform 1 0 444 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1751994658
transform -1 0 556 0 1 105
box -2 -3 98 103
use INVX8  INVX8_4
timestamp 1751994658
transform -1 0 652 0 -1 105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1751994658
transform -1 0 748 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_34
timestamp 1751994658
transform 1 0 556 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1751994658
transform -1 0 612 0 1 105
box -2 -3 34 103
use INVX1  INVX1_74
timestamp 1751994658
transform 1 0 612 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_53
timestamp 1751994658
transform -1 0 676 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_33
timestamp 1751994658
transform -1 0 700 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_32
timestamp 1751994658
transform 1 0 700 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_20
timestamp 1751994658
transform -1 0 756 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1751994658
transform 1 0 748 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_64
timestamp 1751994658
transform 1 0 844 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_33
timestamp 1751994658
transform -1 0 908 0 -1 105
box -2 -3 50 103
use FILL  FILL_0_1_0
timestamp 1751994658
transform -1 0 916 0 -1 105
box -2 -3 10 103
use INVX8  INVX8_6
timestamp 1751994658
transform -1 0 796 0 1 105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1751994658
transform -1 0 892 0 1 105
box -2 -3 98 103
use FILL  FILL_1_1_0
timestamp 1751994658
transform 1 0 892 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1751994658
transform 1 0 900 0 1 105
box -2 -3 10 103
use INVX1  INVX1_80
timestamp 1751994658
transform 1 0 908 0 1 105
box -2 -3 18 103
use FILL  FILL_0_1_1
timestamp 1751994658
transform -1 0 924 0 -1 105
box -2 -3 10 103
use INVX8  INVX8_1
timestamp 1751994658
transform -1 0 964 0 -1 105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1751994658
transform -1 0 1060 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_1
timestamp 1751994658
transform -1 0 1084 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1751994658
transform 1 0 1084 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_65
timestamp 1751994658
transform -1 0 972 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1751994658
transform -1 0 1068 0 1 105
box -2 -3 98 103
use INVX1  INVX1_82
timestamp 1751994658
transform 1 0 1068 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_67
timestamp 1751994658
transform -1 0 1132 0 1 105
box -2 -3 50 103
use INVX8  INVX8_7
timestamp 1751994658
transform -1 0 1220 0 -1 105
box -2 -3 42 103
use NOR2X1  NOR2X1_2
timestamp 1751994658
transform 1 0 1220 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_19
timestamp 1751994658
transform -1 0 1260 0 -1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1751994658
transform 1 0 1260 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_54
timestamp 1751994658
transform 1 0 1132 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_19
timestamp 1751994658
transform 1 0 1148 0 1 105
box -2 -3 50 103
use INVX1  INVX1_83
timestamp 1751994658
transform 1 0 1196 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_68
timestamp 1751994658
transform 1 0 1212 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1751994658
transform 1 0 1260 0 1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_40
timestamp 1751994658
transform -1 0 1420 0 1 105
box -2 -3 50 103
use INVX1  INVX1_53
timestamp 1751994658
transform 1 0 1356 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_40
timestamp 1751994658
transform 1 0 1356 0 -1 105
box -2 -3 26 103
use FILL  FILL_1_2_1
timestamp 1751994658
transform -1 0 1436 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_0
timestamp 1751994658
transform -1 0 1428 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_31
timestamp 1751994658
transform -1 0 1460 0 -1 105
box -2 -3 50 103
use FILL  FILL_0_2_1
timestamp 1751994658
transform -1 0 1412 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_0
timestamp 1751994658
transform -1 0 1404 0 -1 105
box -2 -3 10 103
use INVX1  INVX1_62
timestamp 1751994658
transform 1 0 1380 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_32
timestamp 1751994658
transform -1 0 1484 0 1 105
box -2 -3 50 103
use MUX2X1  MUX2X1_28
timestamp 1751994658
transform 1 0 1460 0 -1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1751994658
transform 1 0 1508 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1751994658
transform 1 0 1604 0 -1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_39
timestamp 1751994658
transform 1 0 1484 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1751994658
transform 1 0 1532 0 1 105
box -2 -3 98 103
use MUX2X1  MUX2X1_27
timestamp 1751994658
transform 1 0 1628 0 1 105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1751994658
transform 1 0 1700 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_1
timestamp 1751994658
transform -1 0 1804 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_23
timestamp 1751994658
transform 1 0 1676 0 1 105
box -2 -3 26 103
use INVX1  INVX1_58
timestamp 1751994658
transform -1 0 1716 0 1 105
box -2 -3 18 103
use INVX1  INVX1_31
timestamp 1751994658
transform 1 0 1716 0 1 105
box -2 -3 18 103
use INVX1  INVX1_25
timestamp 1751994658
transform -1 0 1748 0 1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_35
timestamp 1751994658
transform -1 0 1796 0 1 105
box -2 -3 50 103
use FILL  FILL_2_1
timestamp 1751994658
transform 1 0 1796 0 1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1751994658
transform 1 0 4 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_78
timestamp 1751994658
transform 1 0 100 0 -1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_57
timestamp 1751994658
transform -1 0 164 0 -1 305
box -2 -3 50 103
use AOI22X1  AOI22X1_20
timestamp 1751994658
transform 1 0 164 0 -1 305
box -2 -3 42 103
use CLKBUF1  CLKBUF1_10
timestamp 1751994658
transform -1 0 276 0 -1 305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1751994658
transform 1 0 276 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_0_0
timestamp 1751994658
transform 1 0 372 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1751994658
transform 1 0 380 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_53
timestamp 1751994658
transform 1 0 388 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_12
timestamp 1751994658
transform -1 0 452 0 -1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_50
timestamp 1751994658
transform -1 0 476 0 -1 305
box -2 -3 26 103
use NAND3X1  NAND3X1_14
timestamp 1751994658
transform -1 0 508 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1751994658
transform 1 0 508 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_3
timestamp 1751994658
transform -1 0 556 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_10
timestamp 1751994658
transform 1 0 556 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_27
timestamp 1751994658
transform -1 0 596 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_8
timestamp 1751994658
transform 1 0 596 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_11
timestamp 1751994658
transform -1 0 644 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_11
timestamp 1751994658
transform -1 0 668 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_26
timestamp 1751994658
transform -1 0 684 0 -1 305
box -2 -3 18 103
use OR2X2  OR2X2_2
timestamp 1751994658
transform -1 0 716 0 -1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_2
timestamp 1751994658
transform -1 0 780 0 -1 305
box -2 -3 66 103
use NAND2X1  NAND2X1_9
timestamp 1751994658
transform 1 0 780 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_24
timestamp 1751994658
transform -1 0 820 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1751994658
transform -1 0 916 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_1_0
timestamp 1751994658
transform 1 0 916 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1751994658
transform 1 0 924 0 -1 305
box -2 -3 10 103
use INVX1  INVX1_81
timestamp 1751994658
transform 1 0 932 0 -1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_66
timestamp 1751994658
transform -1 0 996 0 -1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_64
timestamp 1751994658
transform 1 0 996 0 -1 305
box -2 -3 50 103
use INVX1  INVX1_79
timestamp 1751994658
transform -1 0 1060 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1751994658
transform -1 0 1156 0 -1 305
box -2 -3 98 103
use NAND2X1  NAND2X1_34
timestamp 1751994658
transform -1 0 1180 0 -1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_71
timestamp 1751994658
transform 1 0 1180 0 -1 305
box -2 -3 50 103
use INVX1  INVX1_86
timestamp 1751994658
transform -1 0 1244 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_51
timestamp 1751994658
transform -1 0 1268 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1751994658
transform -1 0 1364 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_12
timestamp 1751994658
transform -1 0 1396 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_2_0
timestamp 1751994658
transform -1 0 1404 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1751994658
transform -1 0 1412 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_46
timestamp 1751994658
transform -1 0 1436 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_63
timestamp 1751994658
transform 1 0 1436 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1751994658
transform -1 0 1548 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_46
timestamp 1751994658
transform 1 0 1548 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_12
timestamp 1751994658
transform -1 0 1588 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_49
timestamp 1751994658
transform -1 0 1604 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1751994658
transform 1 0 1604 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_51
timestamp 1751994658
transform -1 0 1716 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_6
timestamp 1751994658
transform -1 0 1748 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1751994658
transform 1 0 1748 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_18
timestamp 1751994658
transform -1 0 1804 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1751994658
transform 1 0 4 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_95
timestamp 1751994658
transform -1 0 148 0 1 305
box -2 -3 50 103
use AOI22X1  AOI22X1_22
timestamp 1751994658
transform 1 0 148 0 1 305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1751994658
transform 1 0 188 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_56
timestamp 1751994658
transform 1 0 284 0 1 305
box -2 -3 50 103
use INVX1  INVX1_77
timestamp 1751994658
transform -1 0 348 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_51
timestamp 1751994658
transform 1 0 348 0 1 305
box -2 -3 50 103
use FILL  FILL_3_0_0
timestamp 1751994658
transform -1 0 404 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1751994658
transform -1 0 412 0 1 305
box -2 -3 10 103
use INVX1  INVX1_72
timestamp 1751994658
transform -1 0 428 0 1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_27
timestamp 1751994658
transform -1 0 460 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_26
timestamp 1751994658
transform 1 0 460 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1751994658
transform 1 0 492 0 1 305
box -2 -3 34 103
use INVX2  INVX2_4
timestamp 1751994658
transform -1 0 540 0 1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_31
timestamp 1751994658
transform 1 0 540 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1751994658
transform -1 0 596 0 1 305
box -2 -3 26 103
use OR2X2  OR2X2_1
timestamp 1751994658
transform -1 0 628 0 1 305
box -2 -3 34 103
use INVX1  INVX1_23
timestamp 1751994658
transform 1 0 628 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_6
timestamp 1751994658
transform 1 0 644 0 1 305
box -2 -3 26 103
use NOR3X1  NOR3X1_4
timestamp 1751994658
transform 1 0 668 0 1 305
box -2 -3 66 103
use NAND2X1  NAND2X1_5
timestamp 1751994658
transform -1 0 756 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_5
timestamp 1751994658
transform -1 0 780 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_12
timestamp 1751994658
transform 1 0 780 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_8
timestamp 1751994658
transform -1 0 828 0 1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_21
timestamp 1751994658
transform -1 0 868 0 1 305
box -2 -3 42 103
use FILL  FILL_3_1_0
timestamp 1751994658
transform 1 0 868 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1751994658
transform 1 0 876 0 1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_99
timestamp 1751994658
transform 1 0 884 0 1 305
box -2 -3 50 103
use INVX1  INVX1_108
timestamp 1751994658
transform -1 0 948 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1751994658
transform 1 0 948 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_37
timestamp 1751994658
transform 1 0 1044 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_24
timestamp 1751994658
transform -1 0 1100 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1751994658
transform -1 0 1196 0 1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_15
timestamp 1751994658
transform 1 0 1196 0 1 305
box -2 -3 34 103
use OR2X2  OR2X2_3
timestamp 1751994658
transform 1 0 1228 0 1 305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_1
timestamp 1751994658
transform -1 0 1332 0 1 305
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1751994658
transform 1 0 1332 0 1 305
box -2 -3 98 103
use FILL  FILL_3_2_0
timestamp 1751994658
transform -1 0 1436 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1751994658
transform -1 0 1444 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_14
timestamp 1751994658
transform -1 0 1476 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1751994658
transform 1 0 1476 0 1 305
box -2 -3 98 103
use INVX1  INVX1_50
timestamp 1751994658
transform 1 0 1572 0 1 305
box -2 -3 18 103
use INVX1  INVX1_57
timestamp 1751994658
transform 1 0 1588 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_26
timestamp 1751994658
transform -1 0 1652 0 1 305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1751994658
transform -1 0 1748 0 1 305
box -2 -3 98 103
use MUX2X1  MUX2X1_59
timestamp 1751994658
transform 1 0 1748 0 1 305
box -2 -3 50 103
use FILL  FILL_4_1
timestamp 1751994658
transform 1 0 1796 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1751994658
transform 1 0 4 0 -1 505
box -2 -3 98 103
use INVX1  INVX1_104
timestamp 1751994658
transform 1 0 100 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_11
timestamp 1751994658
transform -1 0 164 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_12
timestamp 1751994658
transform -1 0 180 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_55
timestamp 1751994658
transform 1 0 180 0 -1 505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_3
timestamp 1751994658
transform -1 0 276 0 -1 505
box -2 -3 74 103
use MUX2X1  MUX2X1_14
timestamp 1751994658
transform 1 0 276 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_15
timestamp 1751994658
transform -1 0 340 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_0_0
timestamp 1751994658
transform 1 0 340 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1751994658
transform 1 0 348 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1751994658
transform 1 0 356 0 -1 505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_9
timestamp 1751994658
transform 1 0 452 0 -1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_1
timestamp 1751994658
transform 1 0 524 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_18
timestamp 1751994658
transform -1 0 580 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_10
timestamp 1751994658
transform -1 0 604 0 -1 505
box -2 -3 26 103
use NOR3X1  NOR3X1_1
timestamp 1751994658
transform -1 0 668 0 -1 505
box -2 -3 66 103
use NAND2X1  NAND2X1_3
timestamp 1751994658
transform 1 0 668 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1751994658
transform -1 0 708 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1751994658
transform 1 0 708 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1751994658
transform 1 0 804 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_1_0
timestamp 1751994658
transform 1 0 900 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1751994658
transform 1 0 908 0 -1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_96
timestamp 1751994658
transform 1 0 916 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_105
timestamp 1751994658
transform -1 0 980 0 -1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_10
timestamp 1751994658
transform 1 0 980 0 -1 505
box -2 -3 42 103
use AOI22X1  AOI22X1_1
timestamp 1751994658
transform 1 0 1020 0 -1 505
box -2 -3 42 103
use INVX2  INVX2_5
timestamp 1751994658
transform 1 0 1060 0 -1 505
box -2 -3 18 103
use INVX1  INVX1_45
timestamp 1751994658
transform 1 0 1076 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1751994658
transform 1 0 1092 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_10
timestamp 1751994658
transform -1 0 1220 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_56
timestamp 1751994658
transform 1 0 1220 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_16
timestamp 1751994658
transform 1 0 1236 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_49
timestamp 1751994658
transform -1 0 1316 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_48
timestamp 1751994658
transform 1 0 1316 0 -1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_46
timestamp 1751994658
transform 1 0 1332 0 -1 505
box -2 -3 50 103
use INVX1  INVX1_44
timestamp 1751994658
transform -1 0 1396 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_2_0
timestamp 1751994658
transform -1 0 1404 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1751994658
transform -1 0 1412 0 -1 505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_6
timestamp 1751994658
transform -1 0 1484 0 -1 505
box -2 -3 74 103
use MUX2X1  MUX2X1_94
timestamp 1751994658
transform 1 0 1484 0 -1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_2
timestamp 1751994658
transform 1 0 1532 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1751994658
transform -1 0 1660 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_13
timestamp 1751994658
transform 1 0 1660 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1751994658
transform -1 0 1708 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1751994658
transform -1 0 1804 0 -1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_79
timestamp 1751994658
transform -1 0 52 0 1 505
box -2 -3 50 103
use INVX1  INVX1_94
timestamp 1751994658
transform -1 0 68 0 1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_23
timestamp 1751994658
transform -1 0 108 0 1 505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1751994658
transform 1 0 108 0 1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_62
timestamp 1751994658
transform -1 0 228 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_60
timestamp 1751994658
transform 1 0 228 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_10
timestamp 1751994658
transform 1 0 252 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_21
timestamp 1751994658
transform -1 0 308 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1751994658
transform 1 0 308 0 1 505
box -2 -3 98 103
use FILL  FILL_5_0_0
timestamp 1751994658
transform 1 0 404 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1751994658
transform 1 0 412 0 1 505
box -2 -3 10 103
use AOI22X1  AOI22X1_6
timestamp 1751994658
transform 1 0 420 0 1 505
box -2 -3 42 103
use NAND3X1  NAND3X1_8
timestamp 1751994658
transform -1 0 492 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_22
timestamp 1751994658
transform -1 0 516 0 1 505
box -2 -3 26 103
use INVX4  INVX4_2
timestamp 1751994658
transform -1 0 540 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_30
timestamp 1751994658
transform 1 0 540 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1751994658
transform -1 0 660 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_4
timestamp 1751994658
transform -1 0 684 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_7
timestamp 1751994658
transform 1 0 684 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_9
timestamp 1751994658
transform -1 0 732 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_98
timestamp 1751994658
transform 1 0 732 0 1 505
box -2 -3 50 103
use INVX1  INVX1_107
timestamp 1751994658
transform -1 0 796 0 1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_7
timestamp 1751994658
transform 1 0 796 0 1 505
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1751994658
transform -1 0 932 0 1 505
box -2 -3 98 103
use FILL  FILL_5_1_0
timestamp 1751994658
transform 1 0 932 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1751994658
transform 1 0 940 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_33
timestamp 1751994658
transform 1 0 948 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1751994658
transform 1 0 980 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1751994658
transform -1 0 1100 0 1 505
box -2 -3 98 103
use INVX1  INVX1_110
timestamp 1751994658
transform 1 0 1100 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_102
timestamp 1751994658
transform -1 0 1164 0 1 505
box -2 -3 50 103
use INVX1  INVX1_43
timestamp 1751994658
transform 1 0 1164 0 1 505
box -2 -3 18 103
use INVX4  INVX4_4
timestamp 1751994658
transform 1 0 1180 0 1 505
box -2 -3 26 103
use NOR3X1  NOR3X1_18
timestamp 1751994658
transform -1 0 1268 0 1 505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1751994658
transform -1 0 1364 0 1 505
box -2 -3 98 103
use INVX1  INVX1_47
timestamp 1751994658
transform 1 0 1364 0 1 505
box -2 -3 18 103
use FILL  FILL_5_2_0
timestamp 1751994658
transform -1 0 1388 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1751994658
transform -1 0 1396 0 1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_24
timestamp 1751994658
transform -1 0 1444 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1751994658
transform 1 0 1444 0 1 505
box -2 -3 98 103
use MUX2X1  MUX2X1_63
timestamp 1751994658
transform 1 0 1540 0 1 505
box -2 -3 50 103
use NOR3X1  NOR3X1_16
timestamp 1751994658
transform 1 0 1588 0 1 505
box -2 -3 66 103
use MUX2X1  MUX2X1_25
timestamp 1751994658
transform 1 0 1652 0 1 505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1751994658
transform -1 0 1796 0 1 505
box -2 -3 98 103
use FILL  FILL_6_1
timestamp 1751994658
transform 1 0 1796 0 1 505
box -2 -3 10 103
use INVX8  INVX8_8
timestamp 1751994658
transform 1 0 4 0 -1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_76
timestamp 1751994658
transform 1 0 44 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1751994658
transform -1 0 188 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_92
timestamp 1751994658
transform 1 0 188 0 -1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_38
timestamp 1751994658
transform -1 0 260 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_103
timestamp 1751994658
transform -1 0 276 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1751994658
transform -1 0 372 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_0_0
timestamp 1751994658
transform -1 0 380 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1751994658
transform -1 0 388 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1751994658
transform -1 0 484 0 -1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_14
timestamp 1751994658
transform 1 0 484 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_25
timestamp 1751994658
transform 1 0 516 0 -1 705
box -2 -3 26 103
use NOR3X1  NOR3X1_19
timestamp 1751994658
transform 1 0 540 0 -1 705
box -2 -3 66 103
use NOR2X1  NOR2X1_33
timestamp 1751994658
transform 1 0 604 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1751994658
transform -1 0 660 0 -1 705
box -2 -3 34 103
use INVX4  INVX4_3
timestamp 1751994658
transform -1 0 684 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_1
timestamp 1751994658
transform 1 0 684 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1751994658
transform 1 0 700 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_66
timestamp 1751994658
transform 1 0 796 0 -1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_43
timestamp 1751994658
transform -1 0 860 0 -1 705
box -2 -3 50 103
use AOI22X1  AOI22X1_5
timestamp 1751994658
transform -1 0 900 0 -1 705
box -2 -3 42 103
use FILL  FILL_6_1_0
timestamp 1751994658
transform -1 0 908 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1751994658
transform -1 0 916 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1751994658
transform -1 0 1012 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_96
timestamp 1751994658
transform 1 0 1012 0 -1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_81
timestamp 1751994658
transform -1 0 1076 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1751994658
transform 1 0 1076 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_28
timestamp 1751994658
transform 1 0 1172 0 -1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_1
timestamp 1751994658
transform 1 0 1196 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1751994658
transform 1 0 1244 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_1
timestamp 1751994658
transform 1 0 1340 0 -1 705
box -2 -3 18 103
use OAI22X1  OAI22X1_8
timestamp 1751994658
transform -1 0 1396 0 -1 705
box -2 -3 42 103
use FILL  FILL_6_2_0
timestamp 1751994658
transform -1 0 1404 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1751994658
transform -1 0 1412 0 -1 705
box -2 -3 10 103
use OAI22X1  OAI22X1_6
timestamp 1751994658
transform -1 0 1452 0 -1 705
box -2 -3 42 103
use NOR3X1  NOR3X1_14
timestamp 1751994658
transform 1 0 1452 0 -1 705
box -2 -3 66 103
use AOI21X1  AOI21X1_8
timestamp 1751994658
transform 1 0 1516 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1751994658
transform -1 0 1580 0 -1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_93
timestamp 1751994658
transform -1 0 1628 0 -1 705
box -2 -3 50 103
use OAI22X1  OAI22X1_7
timestamp 1751994658
transform -1 0 1668 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_19
timestamp 1751994658
transform -1 0 1692 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1751994658
transform -1 0 1788 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_35
timestamp 1751994658
transform 1 0 1788 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1751994658
transform 1 0 4 0 1 705
box -2 -3 98 103
use INVX1  INVX1_91
timestamp 1751994658
transform -1 0 116 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_39
timestamp 1751994658
transform 1 0 116 0 1 705
box -2 -3 26 103
use INVX1  INVX1_75
timestamp 1751994658
transform 1 0 140 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_54
timestamp 1751994658
transform -1 0 204 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_35
timestamp 1751994658
transform 1 0 204 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_20
timestamp 1751994658
transform 1 0 228 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1751994658
transform 1 0 260 0 1 705
box -2 -3 98 103
use INVX1  INVX1_16
timestamp 1751994658
transform 1 0 356 0 1 705
box -2 -3 18 103
use FILL  FILL_7_0_0
timestamp 1751994658
transform -1 0 380 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1751994658
transform -1 0 388 0 1 705
box -2 -3 10 103
use MUX2X1  MUX2X1_15
timestamp 1751994658
transform -1 0 436 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_45
timestamp 1751994658
transform 1 0 436 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1751994658
transform 1 0 460 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_54
timestamp 1751994658
transform -1 0 580 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1751994658
transform -1 0 676 0 1 705
box -2 -3 98 103
use INVX1  INVX1_102
timestamp 1751994658
transform 1 0 676 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_87
timestamp 1751994658
transform -1 0 740 0 1 705
box -2 -3 50 103
use NAND3X1  NAND3X1_16
timestamp 1751994658
transform -1 0 772 0 1 705
box -2 -3 34 103
use INVX2  INVX2_2
timestamp 1751994658
transform -1 0 788 0 1 705
box -2 -3 18 103
use INVX1  INVX1_106
timestamp 1751994658
transform -1 0 804 0 1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_4
timestamp 1751994658
transform 1 0 804 0 1 705
box -2 -3 42 103
use FILL  FILL_7_1_0
timestamp 1751994658
transform -1 0 852 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1751994658
transform -1 0 860 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1751994658
transform -1 0 956 0 1 705
box -2 -3 98 103
use NAND2X1  NAND2X1_59
timestamp 1751994658
transform 1 0 956 0 1 705
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1751994658
transform -1 0 1004 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_46
timestamp 1751994658
transform -1 0 1028 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_35
timestamp 1751994658
transform 1 0 1028 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_100
timestamp 1751994658
transform 1 0 1052 0 1 705
box -2 -3 50 103
use OAI21X1  OAI21X1_9
timestamp 1751994658
transform 1 0 1100 0 1 705
box -2 -3 34 103
use INVX1  INVX1_42
timestamp 1751994658
transform -1 0 1148 0 1 705
box -2 -3 18 103
use NOR3X1  NOR3X1_12
timestamp 1751994658
transform -1 0 1212 0 1 705
box -2 -3 66 103
use OAI22X1  OAI22X1_5
timestamp 1751994658
transform -1 0 1252 0 1 705
box -2 -3 42 103
use MUX2X1  MUX2X1_38
timestamp 1751994658
transform 1 0 1252 0 1 705
box -2 -3 50 103
use INVX1  INVX1_41
timestamp 1751994658
transform -1 0 1316 0 1 705
box -2 -3 18 103
use MUX2X1  MUX2X1_62
timestamp 1751994658
transform -1 0 1364 0 1 705
box -2 -3 50 103
use FILL  FILL_7_2_0
timestamp 1751994658
transform -1 0 1372 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1751994658
transform -1 0 1380 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1751994658
transform -1 0 1476 0 1 705
box -2 -3 98 103
use DFFSR  DFFSR_8
timestamp 1751994658
transform 1 0 1476 0 1 705
box -2 -3 178 103
use MUX2X1  MUX2X1_89
timestamp 1751994658
transform 1 0 1652 0 1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1751994658
transform -1 0 1796 0 1 705
box -2 -3 98 103
use FILL  FILL_8_1
timestamp 1751994658
transform 1 0 1796 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1751994658
transform 1 0 4 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_32
timestamp 1751994658
transform -1 0 132 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_45
timestamp 1751994658
transform -1 0 156 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_52
timestamp 1751994658
transform 1 0 156 0 -1 905
box -2 -3 26 103
use AND2X2  AND2X2_1
timestamp 1751994658
transform -1 0 212 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_58
timestamp 1751994658
transform 1 0 212 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_18
timestamp 1751994658
transform -1 0 268 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1751994658
transform -1 0 292 0 -1 905
box -2 -3 26 103
use NOR3X1  NOR3X1_13
timestamp 1751994658
transform 1 0 292 0 -1 905
box -2 -3 66 103
use NAND3X1  NAND3X1_30
timestamp 1751994658
transform 1 0 356 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_0_0
timestamp 1751994658
transform -1 0 396 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1751994658
transform -1 0 404 0 -1 905
box -2 -3 10 103
use AOI22X1  AOI22X1_17
timestamp 1751994658
transform -1 0 444 0 -1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_36
timestamp 1751994658
transform 1 0 444 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1751994658
transform -1 0 564 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_17
timestamp 1751994658
transform 1 0 564 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_29
timestamp 1751994658
transform 1 0 596 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_61
timestamp 1751994658
transform 1 0 620 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_28
timestamp 1751994658
transform -1 0 676 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_7
timestamp 1751994658
transform 1 0 676 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_48
timestamp 1751994658
transform 1 0 700 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1751994658
transform -1 0 756 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_97
timestamp 1751994658
transform 1 0 756 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_21
timestamp 1751994658
transform -1 0 828 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_56
timestamp 1751994658
transform 1 0 828 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_84
timestamp 1751994658
transform 1 0 852 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_1_0
timestamp 1751994658
transform -1 0 876 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1751994658
transform -1 0 884 0 -1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_69
timestamp 1751994658
transform -1 0 932 0 -1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_31
timestamp 1751994658
transform 1 0 932 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1751994658
transform -1 0 988 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_18
timestamp 1751994658
transform -1 0 1036 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1751994658
transform 1 0 1036 0 -1 905
box -2 -3 98 103
use INVX1  INVX1_40
timestamp 1751994658
transform 1 0 1132 0 -1 905
box -2 -3 18 103
use AOI21X1  AOI21X1_5
timestamp 1751994658
transform -1 0 1180 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_41
timestamp 1751994658
transform -1 0 1228 0 -1 905
box -2 -3 50 103
use INVX1  INVX1_55
timestamp 1751994658
transform -1 0 1244 0 -1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1751994658
transform 1 0 1244 0 -1 905
box -2 -3 98 103
use AOI21X1  AOI21X1_6
timestamp 1751994658
transform 1 0 1340 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_17
timestamp 1751994658
transform -1 0 1396 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_2_0
timestamp 1751994658
transform 1 0 1396 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1751994658
transform 1 0 1404 0 -1 905
box -2 -3 10 103
use DFFSR  DFFSR_7
timestamp 1751994658
transform 1 0 1412 0 -1 905
box -2 -3 178 103
use AOI21X1  AOI21X1_7
timestamp 1751994658
transform 1 0 1588 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1751994658
transform -1 0 1644 0 -1 905
box -2 -3 26 103
use OAI22X1  OAI22X1_2
timestamp 1751994658
transform 1 0 1644 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_3
timestamp 1751994658
transform 1 0 1684 0 -1 905
box -2 -3 34 103
use NOR3X1  NOR3X1_6
timestamp 1751994658
transform 1 0 1716 0 -1 905
box -2 -3 66 103
use BUFX2  BUFX2_7
timestamp 1751994658
transform 1 0 1780 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1751994658
transform 1 0 4 0 1 905
box -2 -3 98 103
use INVX1  INVX1_10
timestamp 1751994658
transform 1 0 100 0 1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_9
timestamp 1751994658
transform -1 0 164 0 1 905
box -2 -3 50 103
use AOI22X1  AOI22X1_14
timestamp 1751994658
transform 1 0 164 0 1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_42
timestamp 1751994658
transform -1 0 228 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_29
timestamp 1751994658
transform -1 0 260 0 1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1751994658
transform -1 0 356 0 1 905
box -2 -3 98 103
use NAND3X1  NAND3X1_29
timestamp 1751994658
transform 1 0 356 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1751994658
transform 1 0 388 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1751994658
transform 1 0 396 0 1 905
box -2 -3 10 103
use AND2X2  AND2X2_2
timestamp 1751994658
transform 1 0 404 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_23
timestamp 1751994658
transform -1 0 468 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1751994658
transform 1 0 468 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_17
timestamp 1751994658
transform -1 0 524 0 1 905
box -2 -3 26 103
use NOR3X1  NOR3X1_17
timestamp 1751994658
transform -1 0 588 0 1 905
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1751994658
transform 1 0 588 0 1 905
box -2 -3 98 103
use INVX1  INVX1_109
timestamp 1751994658
transform 1 0 684 0 1 905
box -2 -3 18 103
use MUX2X1  MUX2X1_101
timestamp 1751994658
transform -1 0 748 0 1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1751994658
transform -1 0 844 0 1 905
box -2 -3 98 103
use FILL  FILL_9_1_0
timestamp 1751994658
transform -1 0 852 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1751994658
transform -1 0 860 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1751994658
transform -1 0 956 0 1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_57
timestamp 1751994658
transform 1 0 956 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_2
timestamp 1751994658
transform 1 0 980 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1751994658
transform -1 0 1100 0 1 905
box -2 -3 98 103
use MUX2X1  MUX2X1_70
timestamp 1751994658
transform -1 0 1148 0 1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_16
timestamp 1751994658
transform -1 0 1172 0 1 905
box -2 -3 26 103
use DFFSR  DFFSR_5
timestamp 1751994658
transform -1 0 1348 0 1 905
box -2 -3 178 103
use FILL  FILL_9_2_0
timestamp 1751994658
transform 1 0 1348 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1751994658
transform 1 0 1356 0 1 905
box -2 -3 10 103
use DFFSR  DFFSR_6
timestamp 1751994658
transform 1 0 1364 0 1 905
box -2 -3 178 103
use MUX2X1  MUX2X1_37
timestamp 1751994658
transform -1 0 1588 0 1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_22
timestamp 1751994658
transform -1 0 1636 0 1 905
box -2 -3 50 103
use INVX1  INVX1_33
timestamp 1751994658
transform -1 0 1652 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1751994658
transform -1 0 1748 0 1 905
box -2 -3 98 103
use BUFX2  BUFX2_5
timestamp 1751994658
transform 1 0 1748 0 1 905
box -2 -3 26 103
use BUFX2  BUFX2_6
timestamp 1751994658
transform 1 0 1772 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1751994658
transform 1 0 1796 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1751994658
transform 1 0 4 0 -1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_13
timestamp 1751994658
transform 1 0 100 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_24
timestamp 1751994658
transform -1 0 156 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1751994658
transform 1 0 156 0 -1 1105
box -2 -3 98 103
use AOI22X1  AOI22X1_3
timestamp 1751994658
transform 1 0 252 0 -1 1105
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1751994658
transform 1 0 292 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_0_0
timestamp 1751994658
transform 1 0 388 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1751994658
transform 1 0 396 0 -1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_12
timestamp 1751994658
transform 1 0 404 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_13
timestamp 1751994658
transform -1 0 468 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_16
timestamp 1751994658
transform 1 0 468 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_4
timestamp 1751994658
transform -1 0 524 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_9
timestamp 1751994658
transform -1 0 564 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_22
timestamp 1751994658
transform -1 0 588 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_11
timestamp 1751994658
transform -1 0 620 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_19
timestamp 1751994658
transform 1 0 620 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_37
timestamp 1751994658
transform -1 0 676 0 -1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1751994658
transform -1 0 772 0 -1 1105
box -2 -3 98 103
use NOR3X1  NOR3X1_7
timestamp 1751994658
transform 1 0 772 0 -1 1105
box -2 -3 66 103
use AOI22X1  AOI22X1_15
timestamp 1751994658
transform 1 0 836 0 -1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_28
timestamp 1751994658
transform -1 0 900 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_1_0
timestamp 1751994658
transform -1 0 908 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1751994658
transform -1 0 916 0 -1 1105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_7
timestamp 1751994658
transform -1 0 988 0 -1 1105
box -2 -3 74 103
use AOI22X1  AOI22X1_13
timestamp 1751994658
transform 1 0 988 0 -1 1105
box -2 -3 42 103
use INVX4  INVX4_5
timestamp 1751994658
transform 1 0 1028 0 -1 1105
box -2 -3 26 103
use AOI22X1  AOI22X1_18
timestamp 1751994658
transform 1 0 1052 0 -1 1105
box -2 -3 42 103
use INVX1  INVX1_85
timestamp 1751994658
transform 1 0 1092 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1751994658
transform -1 0 1204 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1751994658
transform 1 0 1204 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1751994658
transform 1 0 1300 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_2_0
timestamp 1751994658
transform 1 0 1396 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1751994658
transform 1 0 1404 0 -1 1105
box -2 -3 10 103
use INVX1  INVX1_29
timestamp 1751994658
transform 1 0 1412 0 -1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_21
timestamp 1751994658
transform -1 0 1476 0 -1 1105
box -2 -3 50 103
use INVX1  INVX1_39
timestamp 1751994658
transform 1 0 1476 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1751994658
transform -1 0 1588 0 -1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_8
timestamp 1751994658
transform 1 0 1588 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_3
timestamp 1751994658
transform 1 0 1620 0 -1 1105
box -2 -3 42 103
use AOI21X1  AOI21X1_2
timestamp 1751994658
transform 1 0 1660 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_34
timestamp 1751994658
transform -1 0 1708 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1751994658
transform -1 0 1804 0 -1 1105
box -2 -3 98 103
use MUX2X1  MUX2X1_72
timestamp 1751994658
transform -1 0 52 0 1 1105
box -2 -3 50 103
use INVX1  INVX1_87
timestamp 1751994658
transform -1 0 68 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1751994658
transform 1 0 68 0 1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_9
timestamp 1751994658
transform 1 0 164 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_20
timestamp 1751994658
transform -1 0 220 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1751994658
transform 1 0 220 0 1 1105
box -2 -3 98 103
use AOI21X1  AOI21X1_25
timestamp 1751994658
transform 1 0 316 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_38
timestamp 1751994658
transform -1 0 372 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_0_0
timestamp 1751994658
transform 1 0 372 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1751994658
transform 1 0 380 0 1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_14
timestamp 1751994658
transform 1 0 388 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_8
timestamp 1751994658
transform 1 0 412 0 1 1105
box -2 -3 50 103
use INVX1  INVX1_9
timestamp 1751994658
transform -1 0 476 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1751994658
transform 1 0 476 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1751994658
transform -1 0 668 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_99
timestamp 1751994658
transform 1 0 668 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_84
timestamp 1751994658
transform -1 0 732 0 1 1105
box -2 -3 50 103
use NOR3X1  NOR3X1_15
timestamp 1751994658
transform 1 0 732 0 1 1105
box -2 -3 66 103
use NAND3X1  NAND3X1_11
timestamp 1751994658
transform -1 0 828 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_43
timestamp 1751994658
transform -1 0 852 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_48
timestamp 1751994658
transform 1 0 852 0 1 1105
box -2 -3 50 103
use FILL  FILL_11_1_0
timestamp 1751994658
transform -1 0 908 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1751994658
transform -1 0 916 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_70
timestamp 1751994658
transform -1 0 932 0 1 1105
box -2 -3 18 103
use AOI22X1  AOI22X1_19
timestamp 1751994658
transform 1 0 932 0 1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_49
timestamp 1751994658
transform -1 0 996 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1751994658
transform -1 0 1092 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_61
timestamp 1751994658
transform 1 0 1092 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_30
timestamp 1751994658
transform -1 0 1156 0 1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1751994658
transform -1 0 1252 0 1 1105
box -2 -3 98 103
use CLKBUF1  CLKBUF1_4
timestamp 1751994658
transform -1 0 1324 0 1 1105
box -2 -3 74 103
use MUX2X1  MUX2X1_90
timestamp 1751994658
transform 1 0 1324 0 1 1105
box -2 -3 50 103
use INVX1  INVX1_32
timestamp 1751994658
transform -1 0 1388 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_2_0
timestamp 1751994658
transform -1 0 1396 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1751994658
transform -1 0 1404 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1751994658
transform -1 0 1500 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_59
timestamp 1751994658
transform -1 0 1516 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1751994658
transform 1 0 1516 0 1 1105
box -2 -3 98 103
use MUX2X1  MUX2X1_29
timestamp 1751994658
transform 1 0 1612 0 1 1105
box -2 -3 50 103
use INVX1  INVX1_60
timestamp 1751994658
transform -1 0 1676 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_29
timestamp 1751994658
transform 1 0 1676 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_5
timestamp 1751994658
transform 1 0 1700 0 1 1105
box -2 -3 34 103
use NOR3X1  NOR3X1_8
timestamp 1751994658
transform 1 0 1732 0 1 1105
box -2 -3 66 103
use FILL  FILL_12_1
timestamp 1751994658
transform 1 0 1796 0 1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_6
timestamp 1751994658
transform -1 0 52 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_7
timestamp 1751994658
transform -1 0 68 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_10
timestamp 1751994658
transform 1 0 68 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_11
timestamp 1751994658
transform -1 0 132 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1751994658
transform 1 0 132 0 -1 1305
box -2 -3 98 103
use NAND3X1  NAND3X1_17
timestamp 1751994658
transform 1 0 228 0 -1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1751994658
transform 1 0 260 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_0_0
timestamp 1751994658
transform 1 0 356 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1751994658
transform 1 0 364 0 -1 1305
box -2 -3 10 103
use MUX2X1  MUX2X1_3
timestamp 1751994658
transform 1 0 372 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_4
timestamp 1751994658
transform -1 0 436 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_50
timestamp 1751994658
transform 1 0 436 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_71
timestamp 1751994658
transform -1 0 500 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1751994658
transform 1 0 500 0 -1 1305
box -2 -3 98 103
use NAND3X1  NAND3X1_3
timestamp 1751994658
transform -1 0 628 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1751994658
transform 1 0 628 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1751994658
transform -1 0 692 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_22
timestamp 1751994658
transform 1 0 692 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1751994658
transform 1 0 724 0 -1 1305
box -2 -3 34 103
use NOR3X1  NOR3X1_5
timestamp 1751994658
transform 1 0 756 0 -1 1305
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1751994658
transform 1 0 820 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_1_0
timestamp 1751994658
transform 1 0 916 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1751994658
transform 1 0 924 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_101
timestamp 1751994658
transform 1 0 932 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_86
timestamp 1751994658
transform -1 0 996 0 -1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_15
timestamp 1751994658
transform -1 0 1020 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1751994658
transform 1 0 1020 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1751994658
transform -1 0 1076 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1751994658
transform -1 0 1172 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1751994658
transform -1 0 1268 0 -1 1305
box -2 -3 98 103
use INVX1  INVX1_97
timestamp 1751994658
transform 1 0 1268 0 -1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_82
timestamp 1751994658
transform 1 0 1284 0 -1 1305
box -2 -3 50 103
use OAI22X1  OAI22X1_1
timestamp 1751994658
transform -1 0 1372 0 -1 1305
box -2 -3 42 103
use INVX1  INVX1_21
timestamp 1751994658
transform -1 0 1388 0 -1 1305
box -2 -3 18 103
use FILL  FILL_12_2_0
timestamp 1751994658
transform 1 0 1388 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1751994658
transform 1 0 1396 0 -1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_3
timestamp 1751994658
transform 1 0 1404 0 -1 1305
box -2 -3 34 103
use NOR3X1  NOR3X1_3
timestamp 1751994658
transform -1 0 1500 0 -1 1305
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1751994658
transform -1 0 1596 0 -1 1305
box -2 -3 98 103
use OAI22X1  OAI22X1_4
timestamp 1751994658
transform -1 0 1636 0 -1 1305
box -2 -3 42 103
use MUX2X1  MUX2X1_23
timestamp 1751994658
transform 1 0 1636 0 -1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_13
timestamp 1751994658
transform -1 0 1708 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1751994658
transform 1 0 1708 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1751994658
transform 1 0 4 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1751994658
transform 1 0 100 0 1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_5
timestamp 1751994658
transform 1 0 196 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_6
timestamp 1751994658
transform -1 0 260 0 1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_12
timestamp 1751994658
transform 1 0 260 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1751994658
transform 1 0 292 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_9
timestamp 1751994658
transform 1 0 316 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1751994658
transform 1 0 348 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_0_0
timestamp 1751994658
transform 1 0 380 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1751994658
transform 1 0 388 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1751994658
transform 1 0 396 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_39
timestamp 1751994658
transform -1 0 516 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_26
timestamp 1751994658
transform -1 0 548 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_24
timestamp 1751994658
transform 1 0 548 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1751994658
transform 1 0 580 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_2
timestamp 1751994658
transform 1 0 604 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_19
timestamp 1751994658
transform 1 0 636 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_41
timestamp 1751994658
transform -1 0 684 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_42
timestamp 1751994658
transform 1 0 684 0 1 1305
box -2 -3 26 103
use INVX1  INVX1_76
timestamp 1751994658
transform -1 0 724 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_55
timestamp 1751994658
transform 1 0 724 0 1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_20
timestamp 1751994658
transform -1 0 796 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_27
timestamp 1751994658
transform -1 0 820 0 1 1305
box -2 -3 26 103
use NOR3X1  NOR3X1_9
timestamp 1751994658
transform 1 0 820 0 1 1305
box -2 -3 66 103
use FILL  FILL_13_1_0
timestamp 1751994658
transform 1 0 884 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1751994658
transform 1 0 892 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_26
timestamp 1751994658
transform 1 0 900 0 1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_16
timestamp 1751994658
transform 1 0 924 0 1 1305
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1751994658
transform -1 0 1060 0 1 1305
box -2 -3 98 103
use AOI22X1  AOI22X1_8
timestamp 1751994658
transform 1 0 1060 0 1 1305
box -2 -3 42 103
use INVX1  INVX1_67
timestamp 1751994658
transform 1 0 1100 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_44
timestamp 1751994658
transform -1 0 1164 0 1 1305
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1751994658
transform 1 0 1164 0 1 1305
box -2 -3 98 103
use INVX1  INVX1_38
timestamp 1751994658
transform 1 0 1260 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_61
timestamp 1751994658
transform -1 0 1324 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_20
timestamp 1751994658
transform -1 0 1372 0 1 1305
box -2 -3 50 103
use FILL  FILL_13_2_0
timestamp 1751994658
transform -1 0 1380 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1751994658
transform -1 0 1388 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1751994658
transform -1 0 1484 0 1 1305
box -2 -3 98 103
use OAI21X1  OAI21X1_1
timestamp 1751994658
transform -1 0 1516 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_20
timestamp 1751994658
transform 1 0 1516 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_88
timestamp 1751994658
transform -1 0 1580 0 1 1305
box -2 -3 50 103
use NOR3X1  NOR3X1_10
timestamp 1751994658
transform 1 0 1580 0 1 1305
box -2 -3 66 103
use OAI21X1  OAI21X1_7
timestamp 1751994658
transform -1 0 1676 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_34
timestamp 1751994658
transform 1 0 1676 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_91
timestamp 1751994658
transform 1 0 1724 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_36
timestamp 1751994658
transform -1 0 1788 0 1 1305
box -2 -3 18 103
use INVX1  INVX1_28
timestamp 1751994658
transform -1 0 1804 0 1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1751994658
transform 1 0 4 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_41
timestamp 1751994658
transform 1 0 100 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_28
timestamp 1751994658
transform -1 0 156 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1751994658
transform 1 0 156 0 -1 1505
box -2 -3 26 103
use NAND3X1  NAND3X1_13
timestamp 1751994658
transform 1 0 180 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_52
timestamp 1751994658
transform 1 0 212 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_73
timestamp 1751994658
transform -1 0 276 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1751994658
transform -1 0 372 0 -1 1505
box -2 -3 98 103
use FILL  FILL_14_0_0
timestamp 1751994658
transform 1 0 372 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1751994658
transform 1 0 380 0 -1 1505
box -2 -3 10 103
use AOI21X1  AOI21X1_31
timestamp 1751994658
transform 1 0 388 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_44
timestamp 1751994658
transform -1 0 444 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_44
timestamp 1751994658
transform 1 0 444 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1751994658
transform 1 0 468 0 -1 1505
box -2 -3 98 103
use NAND3X1  NAND3X1_25
timestamp 1751994658
transform -1 0 596 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1751994658
transform 1 0 596 0 -1 1505
box -2 -3 26 103
use NOR3X1  NOR3X1_11
timestamp 1751994658
transform 1 0 620 0 -1 1505
box -2 -3 66 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1751994658
transform -1 0 780 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_40
timestamp 1751994658
transform -1 0 804 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_73
timestamp 1751994658
transform 1 0 804 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_88
timestamp 1751994658
transform -1 0 868 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_1_0
timestamp 1751994658
transform -1 0 876 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1751994658
transform -1 0 884 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1751994658
transform -1 0 980 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_32
timestamp 1751994658
transform -1 0 1004 0 -1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_11
timestamp 1751994658
transform -1 0 1044 0 -1 1505
box -2 -3 42 103
use AOI22X1  AOI22X1_2
timestamp 1751994658
transform 1 0 1044 0 -1 1505
box -2 -3 42 103
use INVX1  INVX1_65
timestamp 1751994658
transform 1 0 1084 0 -1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_42
timestamp 1751994658
transform -1 0 1148 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_85
timestamp 1751994658
transform 1 0 1148 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_100
timestamp 1751994658
transform -1 0 1212 0 -1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1751994658
transform -1 0 1308 0 -1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_58
timestamp 1751994658
transform -1 0 1356 0 -1 1505
box -2 -3 50 103
use INVX1  INVX1_22
timestamp 1751994658
transform -1 0 1372 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_2_0
timestamp 1751994658
transform -1 0 1380 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1751994658
transform -1 0 1388 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1751994658
transform -1 0 1484 0 -1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_1
timestamp 1751994658
transform 1 0 1484 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_3
timestamp 1751994658
transform 1 0 1516 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_14
timestamp 1751994658
transform -1 0 1564 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1751994658
transform 1 0 1564 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_15
timestamp 1751994658
transform -1 0 1620 0 -1 1505
box -2 -3 26 103
use DFFSR  DFFSR_2
timestamp 1751994658
transform 1 0 1620 0 -1 1505
box -2 -3 178 103
use FILL  FILL_15_1
timestamp 1751994658
transform -1 0 1804 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1751994658
transform 1 0 4 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_90
timestamp 1751994658
transform 1 0 100 0 1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_75
timestamp 1751994658
transform -1 0 164 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_31
timestamp 1751994658
transform 1 0 164 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_5
timestamp 1751994658
transform -1 0 20 0 -1 1705
box -2 -3 18 103
use MUX2X1  MUX2X1_4
timestamp 1751994658
transform -1 0 68 0 -1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1751994658
transform 1 0 68 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1751994658
transform 1 0 164 0 -1 1705
box -2 -3 98 103
use NAND2X1  NAND2X1_25
timestamp 1751994658
transform 1 0 252 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_89
timestamp 1751994658
transform -1 0 252 0 1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_74
timestamp 1751994658
transform 1 0 188 0 1 1505
box -2 -3 50 103
use FILL  FILL_16_0_1
timestamp 1751994658
transform 1 0 364 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_0
timestamp 1751994658
transform 1 0 356 0 -1 1705
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1751994658
transform 1 0 356 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_0
timestamp 1751994658
transform 1 0 348 0 1 1505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_2
timestamp 1751994658
transform -1 0 348 0 1 1505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1751994658
transform -1 0 356 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1751994658
transform 1 0 364 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_43
timestamp 1751994658
transform 1 0 460 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_30
timestamp 1751994658
transform -1 0 516 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_78
timestamp 1751994658
transform 1 0 516 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_2
timestamp 1751994658
transform 1 0 372 0 -1 1705
box -2 -3 50 103
use INVX1  INVX1_3
timestamp 1751994658
transform -1 0 436 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1751994658
transform 1 0 436 0 -1 1705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_8
timestamp 1751994658
transform -1 0 604 0 -1 1705
box -2 -3 74 103
use INVX1  INVX1_93
timestamp 1751994658
transform -1 0 580 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_48
timestamp 1751994658
transform 1 0 580 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_7
timestamp 1751994658
transform 1 0 604 0 1 1505
box -2 -3 50 103
use INVX1  INVX1_8
timestamp 1751994658
transform -1 0 668 0 1 1505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1751994658
transform -1 0 764 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1751994658
transform 1 0 604 0 -1 1705
box -2 -3 98 103
use INVX8  INVX8_5
timestamp 1751994658
transform 1 0 700 0 -1 1705
box -2 -3 42 103
use INVX8  INVX8_3
timestamp 1751994658
transform 1 0 812 0 -1 1705
box -2 -3 42 103
use CLKBUF1  CLKBUF1_5
timestamp 1751994658
transform 1 0 740 0 -1 1705
box -2 -3 74 103
use AOI21X1  AOI21X1_27
timestamp 1751994658
transform 1 0 764 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1_1
timestamp 1751994658
transform 1 0 900 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_0
timestamp 1751994658
transform 1 0 892 0 -1 1705
box -2 -3 10 103
use INVX8  INVX8_2
timestamp 1751994658
transform 1 0 852 0 -1 1705
box -2 -3 42 103
use MUX2X1  MUX2X1_77
timestamp 1751994658
transform 1 0 908 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_1_1
timestamp 1751994658
transform 1 0 900 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_0
timestamp 1751994658
transform 1 0 892 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1751994658
transform 1 0 908 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1751994658
transform 1 0 796 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_92
timestamp 1751994658
transform -1 0 972 0 1 1505
box -2 -3 18 103
use INVX1  INVX1_69
timestamp 1751994658
transform 1 0 972 0 1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_47
timestamp 1751994658
transform -1 0 1036 0 1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1751994658
transform -1 0 1132 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_80
timestamp 1751994658
transform 1 0 1004 0 -1 1705
box -2 -3 50 103
use INVX1  INVX1_95
timestamp 1751994658
transform -1 0 1068 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1751994658
transform -1 0 1164 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1751994658
transform -1 0 1228 0 1 1505
box -2 -3 98 103
use INVX1  INVX1_68
timestamp 1751994658
transform 1 0 1228 0 1 1505
box -2 -3 18 103
use MUX2X1  MUX2X1_45
timestamp 1751994658
transform -1 0 1292 0 1 1505
box -2 -3 50 103
use DFFSR  DFFSR_3
timestamp 1751994658
transform -1 0 1340 0 -1 1705
box -2 -3 178 103
use MUX2X1  MUX2X1_83
timestamp 1751994658
transform 1 0 1292 0 1 1505
box -2 -3 50 103
use INVX1  INVX1_98
timestamp 1751994658
transform -1 0 1356 0 1 1505
box -2 -3 18 103
use FILL  FILL_15_2_0
timestamp 1751994658
transform 1 0 1356 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1751994658
transform 1 0 1364 0 1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1751994658
transform 1 0 1372 0 1 1505
box -2 -3 98 103
use FILL  FILL_16_2_0
timestamp 1751994658
transform 1 0 1340 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1751994658
transform 1 0 1348 0 -1 1705
box -2 -3 10 103
use DFFSR  DFFSR_1
timestamp 1751994658
transform 1 0 1356 0 -1 1705
box -2 -3 178 103
use CLKBUF1  CLKBUF1_11
timestamp 1751994658
transform 1 0 1468 0 1 1505
box -2 -3 74 103
use INVX1  INVX1_52
timestamp 1751994658
transform 1 0 1540 0 1 1505
box -2 -3 18 103
use DFFSR  DFFSR_4
timestamp 1751994658
transform 1 0 1556 0 1 1505
box -2 -3 178 103
use BUFX2  BUFX2_1
timestamp 1751994658
transform 1 0 1532 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1751994658
transform 1 0 1556 0 -1 1705
box -2 -3 98 103
use BUFX2  BUFX2_3
timestamp 1751994658
transform 1 0 1732 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_30
timestamp 1751994658
transform -1 0 1772 0 1 1505
box -2 -3 18 103
use BUFX2  BUFX2_4
timestamp 1751994658
transform 1 0 1772 0 1 1505
box -2 -3 26 103
use FILL  FILL_16_1
timestamp 1751994658
transform 1 0 1796 0 1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_36
timestamp 1751994658
transform 1 0 1652 0 -1 1705
box -2 -3 50 103
use MUX2X1  MUX2X1_60
timestamp 1751994658
transform 1 0 1700 0 -1 1705
box -2 -3 50 103
use BUFX2  BUFX2_2
timestamp 1751994658
transform 1 0 1748 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1751994658
transform 1 0 1772 0 -1 1705
box -2 -3 26 103
use FILL  FILL_17_1
timestamp 1751994658
transform -1 0 1804 0 -1 1705
box -2 -3 10 103
<< labels >>
flabel metal6 s 368 -30 384 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 888 -30 904 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 598 1728 602 1732 3 FreeSans 24 90 0 0 clk
port 2 nsew
flabel metal2 s 1302 1728 1306 1732 3 FreeSans 24 90 0 0 rst_n
port 3 nsew
flabel metal2 s 1070 -22 1074 -18 7 FreeSans 24 270 0 0 cs
port 4 nsew
flabel metal2 s 1246 -22 1250 -18 7 FreeSans 24 270 0 0 re
port 5 nsew
flabel metal2 s 1086 -22 1090 -18 7 FreeSans 24 270 0 0 we
port 6 nsew
flabel metal2 s 806 -22 810 -18 7 FreeSans 24 270 0 0 addr[0]
port 7 nsew
flabel metal2 s 702 -22 706 -18 7 FreeSans 24 270 0 0 addr[1]
port 8 nsew
flabel metal2 s 614 -22 618 -18 7 FreeSans 24 270 0 0 addr[2]
port 9 nsew
flabel metal2 s 566 -22 570 -18 7 FreeSans 24 270 0 0 addr[3]
port 10 nsew
flabel metal2 s 870 1728 874 1732 3 FreeSans 24 90 0 0 din[0]
port 11 nsew
flabel metal2 s 830 1728 834 1732 3 FreeSans 24 90 0 0 din[1]
port 12 nsew
flabel metal2 s 630 -22 634 -18 7 FreeSans 24 270 0 0 din[2]
port 13 nsew
flabel metal2 s 718 1728 722 1732 3 FreeSans 24 90 0 0 din[3]
port 14 nsew
flabel metal2 s 774 -22 778 -18 7 FreeSans 24 270 0 0 din[4]
port 15 nsew
flabel metal2 s 1198 -22 1202 -18 7 FreeSans 24 270 0 0 din[5]
port 16 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 din[6]
port 17 nsew
flabel metal2 s 942 -22 946 -18 7 FreeSans 24 270 0 0 din[7]
port 18 nsew
flabel metal3 s 1830 1718 1834 1722 3 FreeSans 24 90 0 0 dout[0]
port 19 nsew
flabel metal3 s 1830 1698 1834 1702 3 FreeSans 24 90 0 0 dout[1]
port 20 nsew
flabel metal3 s 1830 1678 1834 1682 3 FreeSans 24 90 0 0 dout[2]
port 21 nsew
flabel metal3 s 1830 1658 1834 1662 3 FreeSans 24 90 0 0 dout[3]
port 22 nsew
flabel metal3 s 1830 1638 1834 1642 3 FreeSans 24 90 0 0 dout[4]
port 23 nsew
flabel metal3 s 1830 1618 1834 1622 3 FreeSans 24 0 0 0 dout[5]
port 24 nsew
flabel metal3 s 1830 1598 1834 1602 3 FreeSans 24 0 0 0 dout[6]
port 25 nsew
flabel metal3 s 1830 1578 1834 1582 3 FreeSans 24 0 0 0 dout[7]
port 26 nsew
<< end >>
