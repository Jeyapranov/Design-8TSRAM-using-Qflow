VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram8t
  CLASS BLOCK ;
  FOREIGN sram8t ;
  ORIGIN 2.600 3.000 ;
  SIZE 186.000 BY 176.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 118.700 165.400 119.100 165.500 ;
        RECT 150.500 165.400 150.900 165.500 ;
        RECT 118.700 165.100 132.200 165.400 ;
        RECT 1.400 160.800 1.800 163.100 ;
        RECT 2.800 160.800 3.200 165.100 ;
        RECT 5.400 160.800 5.800 164.900 ;
        RECT 7.800 160.800 8.200 165.000 ;
        RECT 10.600 160.800 11.000 163.100 ;
        RECT 12.200 160.800 12.600 163.100 ;
        RECT 15.000 160.800 15.400 165.100 ;
        RECT 17.400 160.800 17.800 165.000 ;
        RECT 20.200 160.800 20.600 163.100 ;
        RECT 21.800 160.800 22.200 163.100 ;
        RECT 24.600 160.800 25.000 165.100 ;
        RECT 27.000 160.800 27.400 165.100 ;
        RECT 29.800 160.800 30.200 163.100 ;
        RECT 31.400 160.800 31.800 163.100 ;
        RECT 34.200 160.800 34.600 165.000 ;
        RECT 38.200 160.800 38.600 164.900 ;
        RECT 40.800 160.800 41.200 165.100 ;
        RECT 43.000 160.800 43.400 163.100 ;
        RECT 44.600 160.800 45.000 165.000 ;
        RECT 47.400 160.800 47.800 163.100 ;
        RECT 49.000 160.800 49.400 163.100 ;
        RECT 51.800 160.800 52.200 165.100 ;
        RECT 53.400 160.800 53.800 165.100 ;
        RECT 55.000 160.800 55.400 165.100 ;
        RECT 56.600 160.800 57.000 165.100 ;
        RECT 58.200 160.800 58.600 165.100 ;
        RECT 59.800 160.800 60.200 165.100 ;
        RECT 61.400 160.800 61.800 165.000 ;
        RECT 64.200 160.800 64.600 163.100 ;
        RECT 65.800 160.800 66.200 163.100 ;
        RECT 68.600 160.800 69.000 165.100 ;
        RECT 70.200 160.800 70.600 165.100 ;
        RECT 71.800 160.800 72.200 165.100 ;
        RECT 73.400 160.800 73.800 165.100 ;
        RECT 74.200 160.800 74.600 165.100 ;
        RECT 75.800 160.800 76.200 165.100 ;
        RECT 77.400 160.800 77.800 165.100 ;
        RECT 79.000 160.800 79.400 165.100 ;
        RECT 80.600 160.800 81.000 165.100 ;
        RECT 81.400 160.800 81.800 165.100 ;
        RECT 83.000 160.800 83.400 165.100 ;
        RECT 84.600 160.800 85.000 165.100 ;
        RECT 85.400 160.800 85.800 165.100 ;
        RECT 87.000 160.800 87.400 165.100 ;
        RECT 88.600 160.800 89.000 165.100 ;
        RECT 91.800 160.800 92.200 165.000 ;
        RECT 94.600 160.800 95.000 163.100 ;
        RECT 96.200 160.800 96.600 163.100 ;
        RECT 99.000 160.800 99.400 165.100 ;
        RECT 101.400 160.800 101.800 164.900 ;
        RECT 104.000 160.800 104.400 165.100 ;
        RECT 106.200 160.800 106.600 163.100 ;
        RECT 107.800 160.800 108.200 165.100 ;
        RECT 130.100 165.000 130.500 165.100 ;
        RECT 110.600 160.800 111.000 163.100 ;
        RECT 112.200 160.800 112.600 163.100 ;
        RECT 115.000 160.800 115.400 165.000 ;
        RECT 131.800 164.800 132.200 165.100 ;
        RECT 137.400 165.100 150.900 165.400 ;
        RECT 137.400 164.800 137.800 165.100 ;
        RECT 139.000 165.000 139.500 165.100 ;
        RECT 116.600 160.800 117.000 163.100 ;
        RECT 118.200 160.800 118.600 163.100 ;
        RECT 119.800 160.800 120.200 163.100 ;
        RECT 121.400 160.800 121.800 163.100 ;
        RECT 125.400 160.800 125.800 163.100 ;
        RECT 127.000 160.800 127.400 163.100 ;
        RECT 130.200 160.800 130.600 163.100 ;
        RECT 131.800 160.800 132.200 163.100 ;
        RECT 133.400 160.800 133.800 163.100 ;
        RECT 135.800 160.800 136.200 163.100 ;
        RECT 137.400 160.800 137.800 163.100 ;
        RECT 139.000 160.800 139.400 163.100 ;
        RECT 142.200 160.800 142.600 163.100 ;
        RECT 143.800 160.800 144.200 163.100 ;
        RECT 147.800 160.800 148.200 163.100 ;
        RECT 149.400 160.800 149.800 163.100 ;
        RECT 151.000 160.800 151.400 163.100 ;
        RECT 152.600 160.800 153.000 163.100 ;
        RECT 154.200 160.800 154.600 164.500 ;
        RECT 156.600 160.800 157.000 165.000 ;
        RECT 159.400 160.800 159.800 163.100 ;
        RECT 161.000 160.800 161.400 163.100 ;
        RECT 163.800 160.800 164.200 165.100 ;
        RECT 166.200 160.800 166.600 164.900 ;
        RECT 168.800 160.800 169.200 165.100 ;
        RECT 171.000 160.800 171.400 164.900 ;
        RECT 173.600 160.800 174.000 165.100 ;
        RECT 175.800 160.800 176.200 164.500 ;
        RECT 178.200 160.800 178.600 164.500 ;
        RECT 0.200 160.200 180.600 160.800 ;
        RECT 1.400 156.000 1.800 160.200 ;
        RECT 4.200 157.900 4.600 160.200 ;
        RECT 5.800 157.900 6.200 160.200 ;
        RECT 8.600 155.900 9.000 160.200 ;
        RECT 10.200 157.900 10.600 160.200 ;
        RECT 12.400 155.900 12.800 160.200 ;
        RECT 15.000 156.100 15.400 160.200 ;
        RECT 16.600 157.900 17.000 160.200 ;
        RECT 18.200 157.900 18.600 160.200 ;
        RECT 19.800 156.100 20.200 160.200 ;
        RECT 22.400 155.900 22.800 160.200 ;
        RECT 24.600 157.900 25.000 160.200 ;
        RECT 25.400 157.900 25.800 160.200 ;
        RECT 27.000 157.900 27.400 160.200 ;
        RECT 27.800 155.900 28.200 160.200 ;
        RECT 29.400 155.900 29.800 160.200 ;
        RECT 31.000 155.900 31.400 160.200 ;
        RECT 32.600 155.900 33.000 160.200 ;
        RECT 34.200 155.900 34.600 160.200 ;
        RECT 37.400 156.000 37.800 160.200 ;
        RECT 40.200 157.900 40.600 160.200 ;
        RECT 41.800 157.900 42.200 160.200 ;
        RECT 44.600 155.900 45.000 160.200 ;
        RECT 46.200 155.900 46.600 160.200 ;
        RECT 50.200 156.500 50.600 160.200 ;
        RECT 52.600 156.100 53.000 160.200 ;
        RECT 55.200 155.900 55.600 160.200 ;
        RECT 57.400 157.900 57.800 160.200 ;
        RECT 58.200 157.900 58.600 160.200 ;
        RECT 59.800 157.900 60.200 160.200 ;
        RECT 61.400 156.100 61.800 160.200 ;
        RECT 64.000 155.900 64.400 160.200 ;
        RECT 66.200 157.900 66.600 160.200 ;
        RECT 67.800 155.900 68.200 160.200 ;
        RECT 70.600 157.900 71.000 160.200 ;
        RECT 72.200 157.900 72.600 160.200 ;
        RECT 75.000 156.000 75.400 160.200 ;
        RECT 77.400 156.500 77.800 160.200 ;
        RECT 80.600 156.000 81.000 160.200 ;
        RECT 83.400 157.900 83.800 160.200 ;
        RECT 85.000 157.900 85.400 160.200 ;
        RECT 87.800 155.900 88.200 160.200 ;
        RECT 91.800 156.100 92.200 160.200 ;
        RECT 94.400 155.900 94.800 160.200 ;
        RECT 96.600 157.900 97.000 160.200 ;
        RECT 97.400 157.900 97.800 160.200 ;
        RECT 99.600 155.900 100.000 160.200 ;
        RECT 102.200 156.100 102.600 160.200 ;
        RECT 104.600 155.900 105.000 160.200 ;
        RECT 107.400 157.900 107.800 160.200 ;
        RECT 109.000 157.900 109.400 160.200 ;
        RECT 111.800 156.000 112.200 160.200 ;
        RECT 114.200 155.900 114.600 160.200 ;
        RECT 117.000 157.900 117.400 160.200 ;
        RECT 118.600 157.900 119.000 160.200 ;
        RECT 121.400 156.000 121.800 160.200 ;
        RECT 123.000 157.900 123.400 160.200 ;
        RECT 125.200 155.900 125.600 160.200 ;
        RECT 127.800 156.100 128.200 160.200 ;
        RECT 130.200 156.100 130.600 160.200 ;
        RECT 132.800 155.900 133.200 160.200 ;
        RECT 135.000 157.900 135.400 160.200 ;
        RECT 138.200 156.000 138.600 160.200 ;
        RECT 141.000 157.900 141.400 160.200 ;
        RECT 142.600 157.900 143.000 160.200 ;
        RECT 145.400 155.900 145.800 160.200 ;
        RECT 147.000 155.900 147.400 160.200 ;
        RECT 148.600 155.900 149.000 160.200 ;
        RECT 150.200 155.900 150.600 160.200 ;
        RECT 151.800 155.900 152.200 160.200 ;
        RECT 153.400 155.900 153.800 160.200 ;
        RECT 154.200 157.900 154.600 160.200 ;
        RECT 155.800 157.900 156.200 160.200 ;
        RECT 157.400 157.900 157.800 160.200 ;
        RECT 159.000 157.900 159.400 160.200 ;
        RECT 162.200 157.900 162.600 160.200 ;
        RECT 163.800 157.900 164.200 160.200 ;
        RECT 167.800 157.900 168.200 160.200 ;
        RECT 169.400 157.900 169.800 160.200 ;
        RECT 171.000 157.900 171.400 160.200 ;
        RECT 172.600 157.900 173.000 160.200 ;
        RECT 174.200 156.500 174.600 160.200 ;
        RECT 176.600 157.900 177.000 160.200 ;
        RECT 178.200 156.500 178.600 160.200 ;
        RECT 157.400 155.900 157.800 156.200 ;
        RECT 159.000 155.900 159.500 156.000 ;
        RECT 157.400 155.600 170.900 155.900 ;
        RECT 170.500 155.500 170.900 155.600 ;
        RECT 176.900 145.400 177.300 145.500 ;
        RECT 163.800 145.100 177.300 145.400 ;
        RECT 1.400 140.800 1.800 145.000 ;
        RECT 4.200 140.800 4.600 143.100 ;
        RECT 5.800 140.800 6.200 143.100 ;
        RECT 8.600 140.800 9.000 145.100 ;
        RECT 10.200 140.800 10.600 145.100 ;
        RECT 14.200 140.800 14.600 144.500 ;
        RECT 15.800 140.800 16.200 143.100 ;
        RECT 17.400 140.800 17.800 143.100 ;
        RECT 18.200 140.800 18.600 143.100 ;
        RECT 19.800 140.800 20.200 142.900 ;
        RECT 22.200 140.800 22.600 144.900 ;
        RECT 24.800 140.800 25.200 145.100 ;
        RECT 27.000 140.800 27.400 143.100 ;
        RECT 28.600 140.800 29.000 145.100 ;
        RECT 31.400 140.800 31.800 143.100 ;
        RECT 33.000 140.800 33.400 143.100 ;
        RECT 35.800 140.800 36.200 145.000 ;
        RECT 39.800 140.800 40.200 144.500 ;
        RECT 43.800 140.800 44.200 145.100 ;
        RECT 44.600 140.800 45.000 143.100 ;
        RECT 46.200 140.800 46.600 143.100 ;
        RECT 47.800 140.800 48.200 145.000 ;
        RECT 50.600 140.800 51.000 143.100 ;
        RECT 52.200 140.800 52.600 143.100 ;
        RECT 55.000 140.800 55.400 145.100 ;
        RECT 57.400 140.800 57.800 142.900 ;
        RECT 59.000 140.800 59.400 143.100 ;
        RECT 59.800 140.800 60.200 143.100 ;
        RECT 61.400 140.800 61.800 143.100 ;
        RECT 63.000 140.800 63.400 144.100 ;
        RECT 69.400 140.800 69.800 145.100 ;
        RECT 72.200 140.800 72.600 143.100 ;
        RECT 73.800 140.800 74.200 143.100 ;
        RECT 76.600 140.800 77.000 145.000 ;
        RECT 79.800 140.800 80.200 145.100 ;
        RECT 81.400 140.800 81.800 144.900 ;
        RECT 84.000 140.800 84.400 145.100 ;
        RECT 86.200 140.800 86.600 143.100 ;
        RECT 89.400 140.800 89.800 145.100 ;
        RECT 92.200 140.800 92.600 143.100 ;
        RECT 93.800 140.800 94.200 143.100 ;
        RECT 96.600 140.800 97.000 145.000 ;
        RECT 98.200 140.800 98.600 143.100 ;
        RECT 99.800 140.800 100.200 143.100 ;
        RECT 103.000 140.800 103.400 144.500 ;
        RECT 105.400 140.800 105.800 144.500 ;
        RECT 108.600 140.800 109.000 143.100 ;
        RECT 110.800 140.800 111.200 145.100 ;
        RECT 113.400 140.800 113.800 144.900 ;
        RECT 115.800 140.800 116.200 144.900 ;
        RECT 118.400 140.800 118.800 145.100 ;
        RECT 120.600 140.800 121.000 143.100 ;
        RECT 122.200 140.800 122.600 145.100 ;
        RECT 125.000 140.800 125.400 143.100 ;
        RECT 126.600 140.800 127.000 143.100 ;
        RECT 129.400 140.800 129.800 145.000 ;
        RECT 131.600 140.800 132.000 145.100 ;
        RECT 134.200 140.800 134.600 144.900 ;
        RECT 136.600 140.800 137.000 143.100 ;
        RECT 139.800 140.800 140.200 145.100 ;
        RECT 142.600 140.800 143.000 143.100 ;
        RECT 144.200 140.800 144.600 143.100 ;
        RECT 147.000 140.800 147.400 145.000 ;
        RECT 149.400 140.800 149.800 144.500 ;
        RECT 151.800 140.800 152.200 145.100 ;
        RECT 155.800 140.800 156.200 145.100 ;
        RECT 157.400 140.800 157.800 144.500 ;
        RECT 161.400 140.800 161.800 145.100 ;
        RECT 163.800 144.800 164.200 145.100 ;
        RECT 165.400 145.000 165.900 145.100 ;
        RECT 162.200 140.800 162.600 143.100 ;
        RECT 163.800 140.800 164.200 143.100 ;
        RECT 165.400 140.800 165.800 143.100 ;
        RECT 168.600 140.800 169.000 143.100 ;
        RECT 170.200 140.800 170.600 143.100 ;
        RECT 174.200 140.800 174.600 143.100 ;
        RECT 175.800 140.800 176.200 143.100 ;
        RECT 177.400 140.800 177.800 143.100 ;
        RECT 179.000 140.800 179.400 143.100 ;
        RECT 0.200 140.200 180.600 140.800 ;
        RECT 1.400 136.000 1.800 140.200 ;
        RECT 4.200 137.900 4.600 140.200 ;
        RECT 5.800 137.900 6.200 140.200 ;
        RECT 8.600 135.900 9.000 140.200 ;
        RECT 11.000 136.000 11.400 140.200 ;
        RECT 13.800 137.900 14.200 140.200 ;
        RECT 15.400 137.900 15.800 140.200 ;
        RECT 18.200 135.900 18.600 140.200 ;
        RECT 20.600 136.100 21.000 140.200 ;
        RECT 23.200 135.900 23.600 140.200 ;
        RECT 25.400 137.900 25.800 140.200 ;
        RECT 26.200 137.900 26.600 140.200 ;
        RECT 27.800 138.100 28.200 140.200 ;
        RECT 29.400 137.900 29.800 140.200 ;
        RECT 31.000 137.900 31.400 140.200 ;
        RECT 31.800 137.900 32.200 140.200 ;
        RECT 33.400 138.100 33.800 140.200 ;
        RECT 35.000 137.900 35.400 140.200 ;
        RECT 36.600 138.100 37.000 140.200 ;
        RECT 40.600 136.000 41.000 140.200 ;
        RECT 43.400 137.900 43.800 140.200 ;
        RECT 45.000 137.900 45.400 140.200 ;
        RECT 47.800 135.900 48.200 140.200 ;
        RECT 51.000 135.900 51.400 140.200 ;
        RECT 53.400 136.500 53.800 140.200 ;
        RECT 55.000 137.900 55.400 140.200 ;
        RECT 56.600 138.100 57.000 140.200 ;
        RECT 58.200 137.900 58.600 140.200 ;
        RECT 59.800 137.900 60.200 140.200 ;
        RECT 60.600 137.900 61.000 140.200 ;
        RECT 62.200 138.100 62.600 140.200 ;
        RECT 63.800 137.900 64.200 140.200 ;
        RECT 65.400 137.900 65.800 140.200 ;
        RECT 66.200 137.900 66.600 140.200 ;
        RECT 67.800 137.900 68.200 140.200 ;
        RECT 68.600 137.900 69.000 140.200 ;
        RECT 70.200 137.900 70.600 140.200 ;
        RECT 71.800 137.900 72.200 140.200 ;
        RECT 73.400 136.100 73.800 140.200 ;
        RECT 76.000 135.900 76.400 140.200 ;
        RECT 77.400 137.900 77.800 140.200 ;
        RECT 79.000 137.900 79.400 140.200 ;
        RECT 79.800 137.900 80.200 140.200 ;
        RECT 81.400 137.900 81.800 140.200 ;
        RECT 83.000 136.900 83.400 140.200 ;
        RECT 90.200 137.900 90.600 140.200 ;
        RECT 91.800 137.900 92.200 140.200 ;
        RECT 93.400 136.500 93.800 140.200 ;
        RECT 97.400 135.900 97.800 140.200 ;
        RECT 100.200 137.900 100.600 140.200 ;
        RECT 101.800 137.900 102.200 140.200 ;
        RECT 104.600 136.000 105.000 140.200 ;
        RECT 107.000 136.500 107.400 140.200 ;
        RECT 110.200 137.900 110.600 140.200 ;
        RECT 112.400 135.900 112.800 140.200 ;
        RECT 115.000 136.100 115.400 140.200 ;
        RECT 117.400 136.000 117.800 140.200 ;
        RECT 120.200 137.900 120.600 140.200 ;
        RECT 121.800 137.900 122.200 140.200 ;
        RECT 124.600 135.900 125.000 140.200 ;
        RECT 126.200 137.900 126.600 140.200 ;
        RECT 128.400 135.900 128.800 140.200 ;
        RECT 131.000 136.100 131.400 140.200 ;
        RECT 133.200 135.900 133.600 140.200 ;
        RECT 135.800 136.100 136.200 140.200 ;
        RECT 139.800 135.900 140.200 140.200 ;
        RECT 142.600 137.900 143.000 140.200 ;
        RECT 144.200 137.900 144.600 140.200 ;
        RECT 147.000 136.000 147.400 140.200 ;
        RECT 148.900 137.900 149.300 140.200 ;
        RECT 151.000 135.900 151.400 140.200 ;
        RECT 151.800 137.900 152.200 140.200 ;
        RECT 154.000 135.900 154.400 140.200 ;
        RECT 156.600 136.100 157.000 140.200 ;
        RECT 159.000 136.900 159.400 140.200 ;
        RECT 164.900 137.900 165.300 140.200 ;
        RECT 167.000 135.900 167.400 140.200 ;
        RECT 168.600 136.100 169.000 140.200 ;
        RECT 171.200 135.900 171.600 140.200 ;
        RECT 173.400 136.100 173.800 140.200 ;
        RECT 176.000 135.900 176.400 140.200 ;
        RECT 178.200 137.900 178.600 140.200 ;
        RECT 179.800 137.900 180.200 140.200 ;
        RECT 1.200 120.800 1.600 125.100 ;
        RECT 3.800 120.800 4.200 124.900 ;
        RECT 6.200 120.800 6.600 123.100 ;
        RECT 7.800 120.800 8.200 124.900 ;
        RECT 10.400 120.800 10.800 125.100 ;
        RECT 12.600 120.800 13.000 123.100 ;
        RECT 14.200 120.800 14.600 125.000 ;
        RECT 17.000 120.800 17.400 123.100 ;
        RECT 18.600 120.800 19.000 123.100 ;
        RECT 21.400 120.800 21.800 125.100 ;
        RECT 23.000 120.800 23.400 123.100 ;
        RECT 24.600 120.800 25.000 122.900 ;
        RECT 27.000 120.800 27.400 125.000 ;
        RECT 29.800 120.800 30.200 123.100 ;
        RECT 31.400 120.800 31.800 123.100 ;
        RECT 34.200 120.800 34.600 125.100 ;
        RECT 38.200 120.800 38.600 124.900 ;
        RECT 40.800 120.800 41.200 125.100 ;
        RECT 43.000 120.800 43.400 123.100 ;
        RECT 44.600 120.800 45.000 124.900 ;
        RECT 47.200 120.800 47.600 125.100 ;
        RECT 49.400 120.800 49.800 123.100 ;
        RECT 51.000 120.800 51.400 125.000 ;
        RECT 53.800 120.800 54.200 123.100 ;
        RECT 55.400 120.800 55.800 123.100 ;
        RECT 58.200 120.800 58.600 125.100 ;
        RECT 60.600 120.800 61.000 122.900 ;
        RECT 62.200 120.800 62.600 123.100 ;
        RECT 63.000 120.800 63.400 123.100 ;
        RECT 64.600 120.800 65.000 122.900 ;
        RECT 67.000 120.800 67.400 122.900 ;
        RECT 68.600 120.800 69.000 123.100 ;
        RECT 69.400 120.800 69.800 123.100 ;
        RECT 71.000 120.800 71.400 122.900 ;
        RECT 72.600 120.800 73.000 123.100 ;
        RECT 74.200 120.800 74.600 122.900 ;
        RECT 76.600 120.800 77.000 124.100 ;
        RECT 83.000 120.800 83.400 125.000 ;
        RECT 85.800 120.800 86.200 123.100 ;
        RECT 87.400 120.800 87.800 123.100 ;
        RECT 90.200 120.800 90.600 125.100 ;
        RECT 93.400 120.800 93.800 123.100 ;
        RECT 95.600 120.800 96.000 125.100 ;
        RECT 98.200 120.800 98.600 124.900 ;
        RECT 99.800 120.800 100.200 123.100 ;
        RECT 101.400 120.800 101.800 123.100 ;
        RECT 103.000 120.800 103.400 124.500 ;
        RECT 107.000 120.800 107.400 125.100 ;
        RECT 108.600 120.800 109.000 125.100 ;
        RECT 111.400 120.800 111.800 123.100 ;
        RECT 113.000 120.800 113.400 123.100 ;
        RECT 115.800 120.800 116.200 125.000 ;
        RECT 118.200 120.800 118.600 125.100 ;
        RECT 121.000 120.800 121.400 123.100 ;
        RECT 122.600 120.800 123.000 123.100 ;
        RECT 125.400 120.800 125.800 125.000 ;
        RECT 127.000 120.800 127.400 123.100 ;
        RECT 129.400 120.800 129.800 124.900 ;
        RECT 132.000 120.800 132.400 125.100 ;
        RECT 133.400 120.800 133.800 125.100 ;
        RECT 136.600 120.800 137.000 125.100 ;
        RECT 138.200 120.800 138.600 123.100 ;
        RECT 141.400 120.800 141.800 124.500 ;
        RECT 148.600 120.800 149.000 124.100 ;
        RECT 151.000 120.800 151.400 125.100 ;
        RECT 153.800 120.800 154.200 123.100 ;
        RECT 155.400 120.800 155.800 123.100 ;
        RECT 158.200 120.800 158.600 125.000 ;
        RECT 159.800 120.800 160.200 125.100 ;
        RECT 163.000 120.800 163.400 125.100 ;
        RECT 164.600 120.800 165.000 124.900 ;
        RECT 167.200 120.800 167.600 125.100 ;
        RECT 170.200 120.800 170.600 125.100 ;
        RECT 171.800 120.800 172.200 125.000 ;
        RECT 174.600 120.800 175.000 123.100 ;
        RECT 176.200 120.800 176.600 123.100 ;
        RECT 179.000 120.800 179.400 125.100 ;
        RECT 0.200 120.200 180.600 120.800 ;
        RECT 1.200 115.900 1.600 120.200 ;
        RECT 3.800 116.100 4.200 120.200 ;
        RECT 6.200 117.900 6.600 120.200 ;
        RECT 7.800 116.000 8.200 120.200 ;
        RECT 10.600 117.900 11.000 120.200 ;
        RECT 12.200 117.900 12.600 120.200 ;
        RECT 15.000 115.900 15.400 120.200 ;
        RECT 17.400 116.500 17.800 120.200 ;
        RECT 21.400 115.900 21.800 120.200 ;
        RECT 23.000 116.000 23.400 120.200 ;
        RECT 25.800 117.900 26.200 120.200 ;
        RECT 27.400 117.900 27.800 120.200 ;
        RECT 30.200 115.900 30.600 120.200 ;
        RECT 32.600 116.500 33.000 120.200 ;
        RECT 36.600 115.900 37.000 120.200 ;
        RECT 39.000 117.900 39.400 120.200 ;
        RECT 40.600 117.900 41.000 120.200 ;
        RECT 42.200 116.100 42.600 120.200 ;
        RECT 44.800 115.900 45.200 120.200 ;
        RECT 47.000 117.900 47.400 120.200 ;
        RECT 48.600 116.000 49.000 120.200 ;
        RECT 51.400 117.900 51.800 120.200 ;
        RECT 53.000 117.900 53.400 120.200 ;
        RECT 55.800 115.900 56.200 120.200 ;
        RECT 58.200 115.900 58.600 120.200 ;
        RECT 61.000 117.900 61.400 120.200 ;
        RECT 62.600 117.900 63.000 120.200 ;
        RECT 65.400 116.000 65.800 120.200 ;
        RECT 67.000 117.900 67.400 120.200 ;
        RECT 69.200 115.900 69.600 120.200 ;
        RECT 71.800 116.100 72.200 120.200 ;
        RECT 74.200 116.900 74.600 120.200 ;
        RECT 80.600 118.100 81.000 120.200 ;
        RECT 82.200 117.900 82.600 120.200 ;
        RECT 83.000 117.900 83.400 120.200 ;
        RECT 84.600 117.900 85.000 120.200 ;
        RECT 86.200 116.100 86.600 120.200 ;
        RECT 88.800 115.900 89.200 120.200 ;
        RECT 92.600 117.900 93.000 120.200 ;
        RECT 94.200 116.500 94.600 120.200 ;
        RECT 97.400 117.900 97.800 120.200 ;
        RECT 99.000 117.900 99.400 120.200 ;
        RECT 100.600 115.900 101.000 120.200 ;
        RECT 103.400 117.900 103.800 120.200 ;
        RECT 105.000 117.900 105.400 120.200 ;
        RECT 107.800 116.000 108.200 120.200 ;
        RECT 109.400 117.900 109.800 120.200 ;
        RECT 111.600 115.900 112.000 120.200 ;
        RECT 114.200 116.100 114.600 120.200 ;
        RECT 116.600 115.900 117.000 120.200 ;
        RECT 119.400 117.900 119.800 120.200 ;
        RECT 121.000 117.900 121.400 120.200 ;
        RECT 123.800 116.000 124.200 120.200 ;
        RECT 125.400 115.900 125.800 120.200 ;
        RECT 127.000 115.900 127.400 120.200 ;
        RECT 128.600 115.900 129.000 120.200 ;
        RECT 130.200 115.900 130.600 120.200 ;
        RECT 131.800 115.900 132.200 120.200 ;
        RECT 133.400 116.100 133.800 120.200 ;
        RECT 136.000 115.900 136.400 120.200 ;
        RECT 138.200 117.900 138.600 120.200 ;
        RECT 141.400 115.900 141.800 120.200 ;
        RECT 144.200 117.900 144.600 120.200 ;
        RECT 145.800 117.900 146.200 120.200 ;
        RECT 148.600 116.000 149.000 120.200 ;
        RECT 151.000 117.900 151.400 120.200 ;
        RECT 152.600 116.000 153.000 120.200 ;
        RECT 155.400 117.900 155.800 120.200 ;
        RECT 157.000 117.900 157.400 120.200 ;
        RECT 159.800 115.900 160.200 120.200 ;
        RECT 162.200 116.100 162.600 120.200 ;
        RECT 164.800 115.900 165.200 120.200 ;
        RECT 167.000 117.900 167.400 120.200 ;
        RECT 167.800 117.900 168.200 120.200 ;
        RECT 169.400 117.900 169.800 120.200 ;
        RECT 170.200 115.900 170.600 120.200 ;
        RECT 172.300 117.900 172.700 120.200 ;
        RECT 174.200 116.900 174.600 120.200 ;
        RECT 1.400 100.800 1.800 105.000 ;
        RECT 4.200 100.800 4.600 103.100 ;
        RECT 5.800 100.800 6.200 103.100 ;
        RECT 8.600 100.800 9.000 105.100 ;
        RECT 11.000 100.800 11.400 104.500 ;
        RECT 15.000 100.800 15.400 105.100 ;
        RECT 16.600 100.800 17.000 105.000 ;
        RECT 19.400 100.800 19.800 103.100 ;
        RECT 21.000 100.800 21.400 103.100 ;
        RECT 23.800 100.800 24.200 105.100 ;
        RECT 26.200 100.800 26.600 104.500 ;
        RECT 30.200 100.800 30.600 105.000 ;
        RECT 33.000 100.800 33.400 103.100 ;
        RECT 34.600 100.800 35.000 103.100 ;
        RECT 37.400 100.800 37.800 105.100 ;
        RECT 41.400 100.800 41.800 104.900 ;
        RECT 44.000 100.800 44.400 105.100 ;
        RECT 46.200 100.800 46.600 103.100 ;
        RECT 47.000 100.800 47.400 103.100 ;
        RECT 48.600 100.800 49.000 103.100 ;
        RECT 50.200 100.800 50.600 102.900 ;
        RECT 51.800 100.800 52.200 103.100 ;
        RECT 55.000 100.800 55.400 104.500 ;
        RECT 58.200 100.800 58.600 105.100 ;
        RECT 60.600 100.800 61.000 104.500 ;
        RECT 62.200 100.800 62.600 103.100 ;
        RECT 63.800 100.800 64.200 102.900 ;
        RECT 65.400 100.800 65.800 103.100 ;
        RECT 67.000 100.800 67.400 103.100 ;
        RECT 68.600 100.800 69.000 105.100 ;
        RECT 71.400 100.800 71.800 103.100 ;
        RECT 73.000 100.800 73.400 103.100 ;
        RECT 75.800 100.800 76.200 105.000 ;
        RECT 78.200 100.800 78.600 104.100 ;
        RECT 84.600 100.800 85.000 104.500 ;
        RECT 87.800 100.800 88.200 103.100 ;
        RECT 89.400 100.800 89.800 103.100 ;
        RECT 91.800 100.800 92.200 105.100 ;
        RECT 93.400 100.800 93.800 105.100 ;
        RECT 95.000 100.800 95.400 105.100 ;
        RECT 96.600 100.800 97.000 105.100 ;
        RECT 98.200 100.800 98.600 105.100 ;
        RECT 99.800 100.800 100.200 104.500 ;
        RECT 103.000 100.800 103.400 105.100 ;
        RECT 104.600 100.800 105.000 105.100 ;
        RECT 106.200 100.800 106.600 104.500 ;
        RECT 109.400 100.800 109.800 103.100 ;
        RECT 111.800 100.800 112.200 105.100 ;
        RECT 114.600 100.800 115.000 103.100 ;
        RECT 116.200 100.800 116.600 103.100 ;
        RECT 119.000 100.800 119.400 105.000 ;
        RECT 121.400 100.800 121.800 105.000 ;
        RECT 124.200 100.800 124.600 103.100 ;
        RECT 125.800 100.800 126.200 103.100 ;
        RECT 128.600 100.800 129.000 105.100 ;
        RECT 131.000 100.800 131.400 105.000 ;
        RECT 133.800 100.800 134.200 103.100 ;
        RECT 135.400 100.800 135.800 103.100 ;
        RECT 138.200 100.800 138.600 105.100 ;
        RECT 141.400 100.800 141.800 103.100 ;
        RECT 143.600 100.800 144.000 105.100 ;
        RECT 146.200 100.800 146.600 104.900 ;
        RECT 147.800 100.800 148.200 103.100 ;
        RECT 150.200 100.800 150.600 105.100 ;
        RECT 153.000 100.800 153.400 103.100 ;
        RECT 154.600 100.800 155.000 103.100 ;
        RECT 157.400 100.800 157.800 105.000 ;
        RECT 159.000 100.800 159.400 105.100 ;
        RECT 161.100 100.800 161.500 103.100 ;
        RECT 162.200 100.800 162.600 105.100 ;
        RECT 165.400 100.800 165.800 105.100 ;
        RECT 167.000 100.800 167.400 104.500 ;
        RECT 170.200 100.800 170.600 103.100 ;
        RECT 171.800 100.800 172.200 105.100 ;
        RECT 174.600 100.800 175.000 103.100 ;
        RECT 176.200 100.800 176.600 103.100 ;
        RECT 179.000 100.800 179.400 105.000 ;
        RECT 0.200 100.200 180.600 100.800 ;
        RECT 1.400 96.000 1.800 100.200 ;
        RECT 4.200 97.900 4.600 100.200 ;
        RECT 5.800 97.900 6.200 100.200 ;
        RECT 8.600 95.900 9.000 100.200 ;
        RECT 10.200 97.900 10.600 100.200 ;
        RECT 12.400 95.900 12.800 100.200 ;
        RECT 15.000 96.100 15.400 100.200 ;
        RECT 17.400 96.500 17.800 100.200 ;
        RECT 22.200 95.900 22.600 100.200 ;
        RECT 24.600 96.500 25.000 100.200 ;
        RECT 27.000 95.900 27.400 100.200 ;
        RECT 29.800 97.900 30.200 100.200 ;
        RECT 31.400 97.900 31.800 100.200 ;
        RECT 34.200 96.000 34.600 100.200 ;
        RECT 35.800 97.900 36.200 100.200 ;
        RECT 37.400 98.100 37.800 100.200 ;
        RECT 40.600 97.900 41.000 100.200 ;
        RECT 42.200 96.100 42.600 100.200 ;
        RECT 44.600 98.100 45.000 100.200 ;
        RECT 46.200 97.900 46.600 100.200 ;
        RECT 47.000 97.900 47.400 100.200 ;
        RECT 48.600 98.100 49.000 100.200 ;
        RECT 50.200 97.900 50.600 100.200 ;
        RECT 51.800 97.900 52.200 100.200 ;
        RECT 57.400 96.900 57.800 100.200 ;
        RECT 59.800 96.000 60.200 100.200 ;
        RECT 62.600 97.900 63.000 100.200 ;
        RECT 64.200 97.900 64.600 100.200 ;
        RECT 67.000 95.900 67.400 100.200 ;
        RECT 68.600 97.900 69.000 100.200 ;
        RECT 70.800 95.900 71.200 100.200 ;
        RECT 73.400 96.100 73.800 100.200 ;
        RECT 75.800 95.900 76.200 100.200 ;
        RECT 78.600 97.900 79.000 100.200 ;
        RECT 80.200 97.900 80.600 100.200 ;
        RECT 83.000 96.000 83.400 100.200 ;
        RECT 87.000 95.900 87.400 100.200 ;
        RECT 89.800 97.900 90.200 100.200 ;
        RECT 91.400 97.900 91.800 100.200 ;
        RECT 94.200 96.000 94.600 100.200 ;
        RECT 95.800 97.900 96.200 100.200 ;
        RECT 97.400 97.900 97.800 100.200 ;
        RECT 98.200 97.900 98.600 100.200 ;
        RECT 99.800 97.900 100.200 100.200 ;
        RECT 101.400 95.900 101.800 100.200 ;
        RECT 104.200 97.900 104.600 100.200 ;
        RECT 105.800 97.900 106.200 100.200 ;
        RECT 108.600 96.000 109.000 100.200 ;
        RECT 110.800 95.900 111.200 100.200 ;
        RECT 113.400 96.100 113.800 100.200 ;
        RECT 116.600 95.900 117.000 100.200 ;
        RECT 117.400 97.900 117.800 100.200 ;
        RECT 119.000 97.900 119.400 100.200 ;
        RECT 120.600 97.900 121.000 100.200 ;
        RECT 122.200 97.900 122.600 100.200 ;
        RECT 126.200 97.900 126.600 100.200 ;
        RECT 127.800 97.900 128.200 100.200 ;
        RECT 131.000 97.900 131.400 100.200 ;
        RECT 132.600 97.900 133.000 100.200 ;
        RECT 134.200 97.900 134.600 100.200 ;
        RECT 136.600 97.900 137.000 100.200 ;
        RECT 138.200 97.900 138.600 100.200 ;
        RECT 139.800 97.900 140.200 100.200 ;
        RECT 143.000 97.900 143.400 100.200 ;
        RECT 144.600 97.900 145.000 100.200 ;
        RECT 148.600 97.900 149.000 100.200 ;
        RECT 150.200 97.900 150.600 100.200 ;
        RECT 151.800 97.900 152.200 100.200 ;
        RECT 153.400 97.900 153.800 100.200 ;
        RECT 130.900 95.900 131.400 96.000 ;
        RECT 132.600 95.900 133.000 96.200 ;
        RECT 119.500 95.600 133.000 95.900 ;
        RECT 138.200 95.900 138.600 96.200 ;
        RECT 139.900 95.900 140.300 96.000 ;
        RECT 154.800 95.900 155.200 100.200 ;
        RECT 157.400 96.100 157.800 100.200 ;
        RECT 159.600 95.900 160.000 100.200 ;
        RECT 162.200 96.100 162.600 100.200 ;
        RECT 164.600 97.900 165.000 100.200 ;
        RECT 166.200 95.900 166.600 100.200 ;
        RECT 169.000 97.900 169.400 100.200 ;
        RECT 170.600 97.900 171.000 100.200 ;
        RECT 173.400 96.000 173.800 100.200 ;
        RECT 175.800 96.500 176.200 100.200 ;
        RECT 178.200 96.500 178.600 100.200 ;
        RECT 138.200 95.600 151.700 95.900 ;
        RECT 119.500 95.500 119.900 95.600 ;
        RECT 151.300 95.500 151.700 95.600 ;
        RECT 156.100 85.400 156.500 85.500 ;
        RECT 143.000 85.100 156.500 85.400 ;
        RECT 1.400 80.800 1.800 85.000 ;
        RECT 4.200 80.800 4.600 83.100 ;
        RECT 5.800 80.800 6.200 83.100 ;
        RECT 8.600 80.800 9.000 85.100 ;
        RECT 11.800 80.800 12.200 84.500 ;
        RECT 15.000 80.800 15.400 85.100 ;
        RECT 15.800 80.800 16.200 83.100 ;
        RECT 17.400 80.800 17.800 83.100 ;
        RECT 19.000 80.800 19.400 84.900 ;
        RECT 20.600 80.800 21.000 83.100 ;
        RECT 21.400 80.800 21.800 83.100 ;
        RECT 23.000 80.800 23.400 83.100 ;
        RECT 24.600 80.800 25.000 82.900 ;
        RECT 26.200 80.800 26.600 83.100 ;
        RECT 27.000 80.800 27.400 83.100 ;
        RECT 28.600 80.800 29.000 83.100 ;
        RECT 30.200 80.800 30.600 84.100 ;
        RECT 35.800 80.800 36.200 83.100 ;
        RECT 37.400 80.800 37.800 82.900 ;
        RECT 43.000 80.800 43.400 84.500 ;
        RECT 44.600 80.800 45.000 83.100 ;
        RECT 46.200 80.800 46.600 83.100 ;
        RECT 47.800 80.800 48.200 85.100 ;
        RECT 50.600 80.800 51.000 83.100 ;
        RECT 52.200 80.800 52.600 83.100 ;
        RECT 55.000 80.800 55.400 85.000 ;
        RECT 57.400 80.800 57.800 84.500 ;
        RECT 59.800 80.800 60.200 85.100 ;
        RECT 62.200 80.800 62.600 83.100 ;
        RECT 63.800 80.800 64.200 83.100 ;
        RECT 65.400 80.800 65.800 82.900 ;
        RECT 67.000 80.800 67.400 83.100 ;
        RECT 67.800 80.800 68.200 83.100 ;
        RECT 69.400 80.800 69.800 83.100 ;
        RECT 70.200 80.800 70.600 85.100 ;
        RECT 74.200 80.800 74.600 84.500 ;
        RECT 76.600 80.800 77.000 84.900 ;
        RECT 79.200 80.800 79.600 85.100 ;
        RECT 80.600 80.800 81.000 83.100 ;
        RECT 82.200 80.800 82.600 83.100 ;
        RECT 83.000 80.800 83.400 83.100 ;
        RECT 84.600 80.800 85.000 83.100 ;
        RECT 85.400 80.800 85.800 83.100 ;
        RECT 89.200 80.800 89.600 85.100 ;
        RECT 91.800 80.800 92.200 84.900 ;
        RECT 93.400 80.800 93.800 85.100 ;
        RECT 97.400 80.800 97.800 84.500 ;
        RECT 99.600 80.800 100.000 85.100 ;
        RECT 102.200 80.800 102.600 84.900 ;
        RECT 104.600 80.800 105.000 85.000 ;
        RECT 107.400 80.800 107.800 83.100 ;
        RECT 109.000 80.800 109.400 83.100 ;
        RECT 111.800 80.800 112.200 85.100 ;
        RECT 113.400 80.800 113.800 83.100 ;
        RECT 116.600 80.800 117.000 84.500 ;
        RECT 118.800 80.800 119.200 85.100 ;
        RECT 121.400 80.800 121.800 84.900 ;
        RECT 123.800 80.800 124.200 83.100 ;
        RECT 125.400 80.800 125.800 85.000 ;
        RECT 128.200 80.800 128.600 83.100 ;
        RECT 129.800 80.800 130.200 83.100 ;
        RECT 132.600 80.800 133.000 85.100 ;
        RECT 135.000 80.800 135.400 84.500 ;
        RECT 139.000 80.800 139.400 85.100 ;
        RECT 143.000 84.800 143.400 85.100 ;
        RECT 144.600 85.000 145.100 85.100 ;
        RECT 141.400 80.800 141.800 83.100 ;
        RECT 143.000 80.800 143.400 83.100 ;
        RECT 144.600 80.800 145.000 83.100 ;
        RECT 147.800 80.800 148.200 83.100 ;
        RECT 149.400 80.800 149.800 83.100 ;
        RECT 153.400 80.800 153.800 83.100 ;
        RECT 155.000 80.800 155.400 83.100 ;
        RECT 156.600 80.800 157.000 83.100 ;
        RECT 158.200 80.800 158.600 83.100 ;
        RECT 159.800 80.800 160.200 84.500 ;
        RECT 163.800 80.800 164.200 85.100 ;
        RECT 164.600 80.800 165.000 85.100 ;
        RECT 167.800 80.800 168.200 85.100 ;
        RECT 168.600 80.800 169.000 85.100 ;
        RECT 170.700 80.800 171.100 83.100 ;
        RECT 172.600 80.800 173.000 84.100 ;
        RECT 179.000 80.800 179.400 84.500 ;
        RECT 0.200 80.200 180.600 80.800 ;
        RECT 1.400 76.000 1.800 80.200 ;
        RECT 4.200 77.900 4.600 80.200 ;
        RECT 5.800 77.900 6.200 80.200 ;
        RECT 8.600 75.900 9.000 80.200 ;
        RECT 11.000 77.900 11.400 80.200 ;
        RECT 11.800 77.900 12.200 80.200 ;
        RECT 13.400 77.900 13.800 80.200 ;
        RECT 14.200 77.900 14.600 80.200 ;
        RECT 16.400 75.900 16.800 80.200 ;
        RECT 19.000 76.100 19.400 80.200 ;
        RECT 20.600 77.900 21.000 80.200 ;
        RECT 22.200 77.900 22.600 80.200 ;
        RECT 23.000 77.900 23.400 80.200 ;
        RECT 24.600 78.100 25.000 80.200 ;
        RECT 27.000 76.000 27.400 80.200 ;
        RECT 29.800 77.900 30.200 80.200 ;
        RECT 31.400 77.900 31.800 80.200 ;
        RECT 34.200 75.900 34.600 80.200 ;
        RECT 35.800 77.900 36.200 80.200 ;
        RECT 39.600 75.900 40.000 80.200 ;
        RECT 42.200 76.100 42.600 80.200 ;
        RECT 43.800 77.900 44.200 80.200 ;
        RECT 45.400 77.900 45.800 80.200 ;
        RECT 47.000 76.000 47.400 80.200 ;
        RECT 49.800 77.900 50.200 80.200 ;
        RECT 51.400 77.900 51.800 80.200 ;
        RECT 54.200 75.900 54.600 80.200 ;
        RECT 55.800 77.900 56.200 80.200 ;
        RECT 57.400 77.900 57.800 80.200 ;
        RECT 59.000 75.900 59.400 80.200 ;
        RECT 61.800 77.900 62.200 80.200 ;
        RECT 63.400 77.900 63.800 80.200 ;
        RECT 66.200 76.000 66.600 80.200 ;
        RECT 67.800 77.900 68.200 80.200 ;
        RECT 70.000 75.900 70.400 80.200 ;
        RECT 72.600 76.100 73.000 80.200 ;
        RECT 75.000 78.100 75.400 80.200 ;
        RECT 76.600 77.900 77.000 80.200 ;
        RECT 78.200 75.900 78.600 80.200 ;
        RECT 79.800 77.900 80.200 80.200 ;
        RECT 81.400 76.500 81.800 80.200 ;
        RECT 87.000 75.900 87.400 80.200 ;
        RECT 89.800 77.900 90.200 80.200 ;
        RECT 91.400 77.900 91.800 80.200 ;
        RECT 94.200 76.000 94.600 80.200 ;
        RECT 95.800 77.900 96.200 80.200 ;
        RECT 97.400 77.900 97.800 80.200 ;
        RECT 98.200 75.900 98.600 80.200 ;
        RECT 99.800 75.900 100.200 80.200 ;
        RECT 102.200 75.900 102.600 80.200 ;
        RECT 103.000 75.900 103.400 80.200 ;
        RECT 106.200 76.100 106.600 80.200 ;
        RECT 108.800 75.900 109.200 80.200 ;
        RECT 110.200 75.900 110.600 80.200 ;
        RECT 112.300 77.900 112.700 80.200 ;
        RECT 114.200 77.900 114.600 80.200 ;
        RECT 119.800 76.900 120.200 80.200 ;
        RECT 121.400 75.900 121.800 80.200 ;
        RECT 124.600 75.900 125.000 80.200 ;
        RECT 126.200 76.100 126.600 80.200 ;
        RECT 128.800 75.900 129.200 80.200 ;
        RECT 131.000 77.900 131.400 80.200 ;
        RECT 132.400 75.900 132.800 80.200 ;
        RECT 135.000 76.100 135.400 80.200 ;
        RECT 139.000 75.900 139.400 80.200 ;
        RECT 141.800 77.900 142.200 80.200 ;
        RECT 143.400 77.900 143.800 80.200 ;
        RECT 146.200 76.000 146.600 80.200 ;
        RECT 147.800 77.900 148.200 80.200 ;
        RECT 149.400 77.900 149.800 80.200 ;
        RECT 151.000 77.900 151.400 80.200 ;
        RECT 154.200 77.900 154.600 80.200 ;
        RECT 155.800 77.900 156.200 80.200 ;
        RECT 159.800 77.900 160.200 80.200 ;
        RECT 161.400 77.900 161.800 80.200 ;
        RECT 163.000 77.900 163.400 80.200 ;
        RECT 164.600 77.900 165.000 80.200 ;
        RECT 149.400 75.900 149.800 76.200 ;
        RECT 166.200 76.100 166.600 80.200 ;
        RECT 151.000 75.900 151.500 76.000 ;
        RECT 168.800 75.900 169.200 80.200 ;
        RECT 171.000 75.900 171.400 80.200 ;
        RECT 173.800 77.900 174.200 80.200 ;
        RECT 175.400 77.900 175.800 80.200 ;
        RECT 178.200 76.000 178.600 80.200 ;
        RECT 149.400 75.600 162.900 75.900 ;
        RECT 162.500 75.500 162.900 75.600 ;
        RECT 0.600 60.800 1.000 65.100 ;
        RECT 2.200 60.800 2.600 65.100 ;
        RECT 3.800 60.800 4.200 65.100 ;
        RECT 5.400 60.800 5.800 64.900 ;
        RECT 8.000 60.800 8.400 65.100 ;
        RECT 10.200 60.800 10.600 65.100 ;
        RECT 13.000 60.800 13.400 63.100 ;
        RECT 14.600 60.800 15.000 63.100 ;
        RECT 17.400 60.800 17.800 65.000 ;
        RECT 19.800 60.800 20.200 64.900 ;
        RECT 22.400 60.800 22.800 65.100 ;
        RECT 23.800 60.800 24.200 63.100 ;
        RECT 25.400 60.800 25.800 63.100 ;
        RECT 27.000 60.800 27.400 63.100 ;
        RECT 28.600 60.800 29.000 65.100 ;
        RECT 31.400 60.800 31.800 63.100 ;
        RECT 33.000 60.800 33.400 63.100 ;
        RECT 35.800 60.800 36.200 65.000 ;
        RECT 39.800 60.800 40.200 65.100 ;
        RECT 42.600 60.800 43.000 63.100 ;
        RECT 44.200 60.800 44.600 63.100 ;
        RECT 47.000 60.800 47.400 65.000 ;
        RECT 49.400 60.800 49.800 64.500 ;
        RECT 51.800 60.800 52.200 65.100 ;
        RECT 55.000 60.800 55.400 64.100 ;
        RECT 60.600 60.800 61.000 65.100 ;
        RECT 64.600 60.800 65.000 64.500 ;
        RECT 66.200 60.800 66.600 65.100 ;
        RECT 67.800 60.800 68.200 65.100 ;
        RECT 68.600 60.800 69.000 65.100 ;
        RECT 71.000 60.800 71.400 65.000 ;
        RECT 73.800 60.800 74.200 63.100 ;
        RECT 75.400 60.800 75.800 63.100 ;
        RECT 78.200 60.800 78.600 65.100 ;
        RECT 79.800 60.800 80.200 63.100 ;
        RECT 82.000 60.800 82.400 65.100 ;
        RECT 84.600 60.800 85.000 64.900 ;
        RECT 88.600 60.800 89.000 64.500 ;
        RECT 92.600 60.800 93.000 65.100 ;
        RECT 95.400 60.800 95.800 63.100 ;
        RECT 97.000 60.800 97.400 63.100 ;
        RECT 99.800 60.800 100.200 65.000 ;
        RECT 101.400 60.800 101.800 63.100 ;
        RECT 103.600 60.800 104.000 65.100 ;
        RECT 106.200 60.800 106.600 64.900 ;
        RECT 108.600 60.800 109.000 65.000 ;
        RECT 111.400 60.800 111.800 63.100 ;
        RECT 113.000 60.800 113.400 63.100 ;
        RECT 115.800 60.800 116.200 65.100 ;
        RECT 117.400 60.800 117.800 65.100 ;
        RECT 120.600 60.800 121.000 64.900 ;
        RECT 123.200 60.800 123.600 65.100 ;
        RECT 125.400 60.800 125.800 65.000 ;
        RECT 128.200 60.800 128.600 63.100 ;
        RECT 129.800 60.800 130.200 63.100 ;
        RECT 132.600 60.800 133.000 65.100 ;
        RECT 134.200 60.800 134.600 63.100 ;
        RECT 135.800 60.800 136.200 65.100 ;
        RECT 139.000 60.800 139.400 65.100 ;
        RECT 141.400 60.800 141.800 65.100 ;
        RECT 144.600 60.800 145.000 65.100 ;
        RECT 146.200 60.800 146.600 64.100 ;
        RECT 152.600 60.800 153.000 64.500 ;
        RECT 155.300 60.800 155.700 63.100 ;
        RECT 157.400 60.800 157.800 65.100 ;
        RECT 158.800 60.800 159.200 65.100 ;
        RECT 161.400 60.800 161.800 64.900 ;
        RECT 163.000 60.800 163.400 65.100 ;
        RECT 166.200 60.800 166.600 65.100 ;
        RECT 168.600 60.800 169.000 65.100 ;
        RECT 170.200 60.800 170.600 65.100 ;
        RECT 173.000 60.800 173.400 63.100 ;
        RECT 174.600 60.800 175.000 63.100 ;
        RECT 177.400 60.800 177.800 65.000 ;
        RECT 179.000 60.800 179.400 63.100 ;
        RECT 0.200 60.200 180.600 60.800 ;
        RECT 1.200 55.900 1.600 60.200 ;
        RECT 3.800 56.100 4.200 60.200 ;
        RECT 6.200 57.900 6.600 60.200 ;
        RECT 9.400 56.500 9.800 60.200 ;
        RECT 11.800 56.000 12.200 60.200 ;
        RECT 14.600 57.900 15.000 60.200 ;
        RECT 16.200 57.900 16.600 60.200 ;
        RECT 19.000 55.900 19.400 60.200 ;
        RECT 20.600 57.900 21.000 60.200 ;
        RECT 22.200 57.900 22.600 60.200 ;
        RECT 23.000 57.900 23.400 60.200 ;
        RECT 24.600 57.900 25.000 60.200 ;
        RECT 26.200 56.500 26.600 60.200 ;
        RECT 30.200 55.900 30.600 60.200 ;
        RECT 31.800 56.000 32.200 60.200 ;
        RECT 34.600 57.900 35.000 60.200 ;
        RECT 36.200 57.900 36.600 60.200 ;
        RECT 39.000 55.900 39.400 60.200 ;
        RECT 43.000 56.500 43.400 60.200 ;
        RECT 47.000 58.100 47.400 60.200 ;
        RECT 48.600 57.900 49.000 60.200 ;
        RECT 49.400 57.900 49.800 60.200 ;
        RECT 51.000 57.900 51.400 60.200 ;
        RECT 51.800 55.900 52.200 60.200 ;
        RECT 53.400 55.900 53.800 60.200 ;
        RECT 54.200 55.900 54.600 60.200 ;
        RECT 57.400 55.900 57.800 60.200 ;
        RECT 60.200 57.900 60.600 60.200 ;
        RECT 61.800 57.900 62.200 60.200 ;
        RECT 64.600 56.000 65.000 60.200 ;
        RECT 67.800 55.900 68.200 60.200 ;
        RECT 68.600 55.900 69.000 60.200 ;
        RECT 72.600 55.900 73.000 60.200 ;
        RECT 74.200 56.100 74.600 60.200 ;
        RECT 76.800 55.900 77.200 60.200 ;
        RECT 79.000 57.900 79.400 60.200 ;
        RECT 80.600 56.500 81.000 60.200 ;
        RECT 84.600 55.900 85.000 60.200 ;
        RECT 87.400 57.900 87.800 60.200 ;
        RECT 89.000 57.900 89.400 60.200 ;
        RECT 91.800 56.000 92.200 60.200 ;
        RECT 95.800 56.500 96.200 60.200 ;
        RECT 98.200 55.900 98.600 60.200 ;
        RECT 101.400 55.900 101.800 60.200 ;
        RECT 104.200 57.900 104.600 60.200 ;
        RECT 105.800 57.900 106.200 60.200 ;
        RECT 108.600 56.000 109.000 60.200 ;
        RECT 110.200 57.900 110.600 60.200 ;
        RECT 112.400 55.900 112.800 60.200 ;
        RECT 115.000 56.100 115.400 60.200 ;
        RECT 116.600 57.900 117.000 60.200 ;
        RECT 118.200 55.900 118.600 60.200 ;
        RECT 119.800 55.900 120.200 60.200 ;
        RECT 125.400 56.900 125.800 60.200 ;
        RECT 127.800 55.900 128.200 60.200 ;
        RECT 130.600 57.900 131.000 60.200 ;
        RECT 132.200 57.900 132.600 60.200 ;
        RECT 135.000 56.000 135.400 60.200 ;
        RECT 136.600 57.900 137.000 60.200 ;
        RECT 140.400 55.900 140.800 60.200 ;
        RECT 143.000 56.100 143.400 60.200 ;
        RECT 145.400 56.000 145.800 60.200 ;
        RECT 148.200 57.900 148.600 60.200 ;
        RECT 149.800 57.900 150.200 60.200 ;
        RECT 152.600 55.900 153.000 60.200 ;
        RECT 155.000 56.100 155.400 60.200 ;
        RECT 157.600 55.900 158.000 60.200 ;
        RECT 159.800 56.900 160.200 60.200 ;
        RECT 166.200 56.100 166.600 60.200 ;
        RECT 168.800 55.900 169.200 60.200 ;
        RECT 171.000 55.900 171.400 60.200 ;
        RECT 173.800 57.900 174.200 60.200 ;
        RECT 175.400 57.900 175.800 60.200 ;
        RECT 178.200 56.000 178.600 60.200 ;
        RECT 1.400 40.800 1.800 45.000 ;
        RECT 4.200 40.800 4.600 43.100 ;
        RECT 5.800 40.800 6.200 43.100 ;
        RECT 8.600 40.800 9.000 45.100 ;
        RECT 10.200 40.800 10.600 43.100 ;
        RECT 12.400 40.800 12.800 45.100 ;
        RECT 15.000 40.800 15.400 44.900 ;
        RECT 17.400 40.800 17.800 43.100 ;
        RECT 18.200 40.800 18.600 43.100 ;
        RECT 19.800 40.800 20.200 43.100 ;
        RECT 20.600 40.800 21.000 45.100 ;
        RECT 22.200 40.800 22.600 45.100 ;
        RECT 23.800 40.800 24.200 45.100 ;
        RECT 25.400 40.800 25.800 45.100 ;
        RECT 27.000 40.800 27.400 45.100 ;
        RECT 28.600 40.800 29.000 44.900 ;
        RECT 31.200 40.800 31.600 45.100 ;
        RECT 33.400 40.800 33.800 43.100 ;
        RECT 36.600 40.800 37.000 45.000 ;
        RECT 39.400 40.800 39.800 43.100 ;
        RECT 41.000 40.800 41.400 43.100 ;
        RECT 43.800 40.800 44.200 45.100 ;
        RECT 45.400 40.800 45.800 45.100 ;
        RECT 47.000 40.800 47.400 45.100 ;
        RECT 48.600 40.800 49.000 45.100 ;
        RECT 50.200 40.800 50.600 45.100 ;
        RECT 51.800 40.800 52.200 45.100 ;
        RECT 52.600 40.800 53.000 45.100 ;
        RECT 56.600 40.800 57.000 44.500 ;
        RECT 59.800 40.800 60.200 45.100 ;
        RECT 65.400 40.800 65.800 44.100 ;
        RECT 67.000 40.800 67.400 43.100 ;
        RECT 68.600 40.800 69.000 43.100 ;
        RECT 70.200 40.800 70.600 43.100 ;
        RECT 71.800 40.800 72.200 45.000 ;
        RECT 74.600 40.800 75.000 43.100 ;
        RECT 76.200 40.800 76.600 43.100 ;
        RECT 79.000 40.800 79.400 45.100 ;
        RECT 81.400 40.800 81.800 45.000 ;
        RECT 84.200 40.800 84.600 43.100 ;
        RECT 85.800 40.800 86.200 43.100 ;
        RECT 88.600 40.800 89.000 45.100 ;
        RECT 92.600 40.800 93.000 44.900 ;
        RECT 95.200 40.800 95.600 45.100 ;
        RECT 97.400 40.800 97.800 43.100 ;
        RECT 99.000 40.800 99.400 44.500 ;
        RECT 103.000 40.800 103.400 44.500 ;
        RECT 106.200 40.800 106.600 45.100 ;
        RECT 107.800 40.800 108.200 43.100 ;
        RECT 110.200 40.800 110.600 45.000 ;
        RECT 113.000 40.800 113.400 43.100 ;
        RECT 114.600 40.800 115.000 43.100 ;
        RECT 117.400 40.800 117.800 45.100 ;
        RECT 119.300 40.800 119.700 43.100 ;
        RECT 121.400 40.800 121.800 45.100 ;
        RECT 122.200 40.800 122.600 43.100 ;
        RECT 123.800 40.800 124.200 45.100 ;
        RECT 125.900 40.800 126.300 43.100 ;
        RECT 127.600 40.800 128.000 45.100 ;
        RECT 130.200 40.800 130.600 44.900 ;
        RECT 131.800 40.800 132.200 43.100 ;
        RECT 134.200 40.800 134.600 44.900 ;
        RECT 136.800 40.800 137.200 45.100 ;
        RECT 139.000 40.800 139.400 43.100 ;
        RECT 141.400 40.800 141.800 45.100 ;
        RECT 143.000 40.800 143.400 45.100 ;
        RECT 144.600 40.800 145.000 45.100 ;
        RECT 146.200 40.800 146.600 45.100 ;
        RECT 147.800 40.800 148.200 45.100 ;
        RECT 149.400 40.800 149.800 44.900 ;
        RECT 152.000 40.800 152.400 45.100 ;
        RECT 153.400 40.800 153.800 45.100 ;
        RECT 155.500 40.800 155.900 43.100 ;
        RECT 157.400 40.800 157.800 45.100 ;
        RECT 160.200 40.800 160.600 43.100 ;
        RECT 161.800 40.800 162.200 43.100 ;
        RECT 164.600 40.800 165.000 45.000 ;
        RECT 166.200 40.800 166.600 45.100 ;
        RECT 168.300 40.800 168.700 43.100 ;
        RECT 170.200 40.800 170.600 43.100 ;
        RECT 171.800 40.800 172.200 45.100 ;
        RECT 174.600 40.800 175.000 43.100 ;
        RECT 176.200 40.800 176.600 43.100 ;
        RECT 179.000 40.800 179.400 45.000 ;
        RECT 0.200 40.200 180.600 40.800 ;
        RECT 1.400 36.000 1.800 40.200 ;
        RECT 4.200 37.900 4.600 40.200 ;
        RECT 5.800 37.900 6.200 40.200 ;
        RECT 8.600 35.900 9.000 40.200 ;
        RECT 10.800 35.900 11.200 40.200 ;
        RECT 13.400 36.100 13.800 40.200 ;
        RECT 15.800 36.500 16.200 40.200 ;
        RECT 19.800 36.000 20.200 40.200 ;
        RECT 22.600 37.900 23.000 40.200 ;
        RECT 24.200 37.900 24.600 40.200 ;
        RECT 27.000 35.900 27.400 40.200 ;
        RECT 29.400 36.100 29.800 40.200 ;
        RECT 32.000 35.900 32.400 40.200 ;
        RECT 34.200 37.900 34.600 40.200 ;
        RECT 35.800 36.100 36.200 40.200 ;
        RECT 38.400 35.900 38.800 40.200 ;
        RECT 42.200 37.900 42.600 40.200 ;
        RECT 43.800 38.100 44.200 40.200 ;
        RECT 45.400 37.900 45.800 40.200 ;
        RECT 46.200 37.900 46.600 40.200 ;
        RECT 47.800 38.100 48.200 40.200 ;
        RECT 49.400 37.900 49.800 40.200 ;
        RECT 51.000 38.100 51.400 40.200 ;
        RECT 53.400 35.900 53.800 40.200 ;
        RECT 54.200 37.900 54.600 40.200 ;
        RECT 55.800 38.100 56.200 40.200 ;
        RECT 59.000 35.900 59.400 40.200 ;
        RECT 60.900 35.900 61.300 40.200 ;
        RECT 63.000 37.900 63.400 40.200 ;
        RECT 64.600 37.900 65.000 40.200 ;
        RECT 66.200 37.900 66.600 40.200 ;
        RECT 67.800 36.900 68.200 40.200 ;
        RECT 73.400 37.900 73.800 40.200 ;
        RECT 75.000 37.900 75.400 40.200 ;
        RECT 77.400 35.900 77.800 40.200 ;
        RECT 78.200 35.900 78.600 40.200 ;
        RECT 82.200 35.900 82.600 40.200 ;
        RECT 85.400 36.500 85.800 40.200 ;
        RECT 89.400 36.100 89.800 40.200 ;
        RECT 92.000 35.900 92.400 40.200 ;
        RECT 94.200 37.900 94.600 40.200 ;
        RECT 95.800 36.000 96.200 40.200 ;
        RECT 98.600 37.900 99.000 40.200 ;
        RECT 100.200 37.900 100.600 40.200 ;
        RECT 103.000 35.900 103.400 40.200 ;
        RECT 104.600 35.900 105.000 40.200 ;
        RECT 108.600 36.500 109.000 40.200 ;
        RECT 111.000 35.900 111.400 40.200 ;
        RECT 113.800 37.900 114.200 40.200 ;
        RECT 115.400 37.900 115.800 40.200 ;
        RECT 118.200 36.000 118.600 40.200 ;
        RECT 119.800 35.900 120.200 40.200 ;
        RECT 121.900 37.900 122.300 40.200 ;
        RECT 124.300 35.900 124.700 40.200 ;
        RECT 126.200 35.900 126.600 40.200 ;
        RECT 127.800 35.900 128.200 40.200 ;
        RECT 129.400 35.900 129.800 40.200 ;
        RECT 131.000 35.900 131.400 40.200 ;
        RECT 132.600 35.900 133.000 40.200 ;
        RECT 134.200 36.000 134.600 40.200 ;
        RECT 137.000 37.900 137.400 40.200 ;
        RECT 138.600 37.900 139.000 40.200 ;
        RECT 141.400 35.900 141.800 40.200 ;
        RECT 144.900 37.900 145.300 40.200 ;
        RECT 147.000 35.900 147.400 40.200 ;
        RECT 148.600 36.000 149.000 40.200 ;
        RECT 151.400 37.900 151.800 40.200 ;
        RECT 153.000 37.900 153.400 40.200 ;
        RECT 155.800 35.900 156.200 40.200 ;
        RECT 157.400 37.900 157.800 40.200 ;
        RECT 159.000 37.900 159.400 40.200 ;
        RECT 161.200 35.900 161.600 40.200 ;
        RECT 163.800 36.100 164.200 40.200 ;
        RECT 166.200 35.900 166.600 40.200 ;
        RECT 169.000 37.900 169.400 40.200 ;
        RECT 170.600 37.900 171.000 40.200 ;
        RECT 173.400 36.000 173.800 40.200 ;
        RECT 175.800 36.100 176.200 40.200 ;
        RECT 178.400 35.900 178.800 40.200 ;
        RECT 1.400 20.800 1.800 25.000 ;
        RECT 4.200 20.800 4.600 23.100 ;
        RECT 5.800 20.800 6.200 23.100 ;
        RECT 8.600 20.800 9.000 25.100 ;
        RECT 10.200 20.800 10.600 23.100 ;
        RECT 12.400 20.800 12.800 25.100 ;
        RECT 15.000 20.800 15.400 24.900 ;
        RECT 17.400 20.800 17.800 24.500 ;
        RECT 20.600 20.800 21.000 25.100 ;
        RECT 22.200 20.800 22.600 25.100 ;
        RECT 23.800 20.800 24.200 25.100 ;
        RECT 25.400 20.800 25.800 25.100 ;
        RECT 27.000 20.800 27.400 25.100 ;
        RECT 28.600 20.800 29.000 25.000 ;
        RECT 31.400 20.800 31.800 23.100 ;
        RECT 33.000 20.800 33.400 23.100 ;
        RECT 35.800 20.800 36.200 25.100 ;
        RECT 39.000 20.800 39.400 23.100 ;
        RECT 40.600 20.800 41.000 23.100 ;
        RECT 43.800 20.800 44.200 24.500 ;
        RECT 45.400 20.800 45.800 23.100 ;
        RECT 47.000 20.800 47.400 23.100 ;
        RECT 48.600 20.800 49.000 22.900 ;
        RECT 50.200 20.800 50.600 23.100 ;
        RECT 51.000 20.800 51.400 23.100 ;
        RECT 52.600 20.800 53.000 22.900 ;
        RECT 55.000 20.800 55.400 25.100 ;
        RECT 55.800 20.800 56.200 23.100 ;
        RECT 57.400 20.800 57.800 23.100 ;
        RECT 59.000 20.800 59.400 23.100 ;
        RECT 59.800 20.800 60.200 23.100 ;
        RECT 61.400 20.800 61.800 23.100 ;
        RECT 63.800 20.800 64.200 25.100 ;
        RECT 64.600 20.800 65.000 23.100 ;
        RECT 66.200 20.800 66.600 23.100 ;
        RECT 67.800 20.800 68.200 23.100 ;
        RECT 69.700 20.800 70.100 25.100 ;
        RECT 76.600 20.800 77.000 24.100 ;
        RECT 78.200 20.800 78.600 23.100 ;
        RECT 79.800 20.800 80.200 23.100 ;
        RECT 81.400 20.800 81.800 23.100 ;
        RECT 83.000 20.800 83.400 25.100 ;
        RECT 85.800 20.800 86.200 23.100 ;
        RECT 87.400 20.800 87.800 23.100 ;
        RECT 90.200 20.800 90.600 25.000 ;
        RECT 93.400 20.800 93.800 23.100 ;
        RECT 95.600 20.800 96.000 25.100 ;
        RECT 98.200 20.800 98.600 24.900 ;
        RECT 100.600 20.800 101.000 24.900 ;
        RECT 103.200 20.800 103.600 25.100 ;
        RECT 105.400 20.800 105.800 23.100 ;
        RECT 107.000 20.800 107.400 25.100 ;
        RECT 109.800 20.800 110.200 23.100 ;
        RECT 111.400 20.800 111.800 23.100 ;
        RECT 114.200 20.800 114.600 25.000 ;
        RECT 115.800 20.800 116.200 23.100 ;
        RECT 117.400 20.800 117.800 23.100 ;
        RECT 119.000 20.800 119.400 24.900 ;
        RECT 121.600 20.800 122.000 25.100 ;
        RECT 123.800 20.800 124.200 23.100 ;
        RECT 124.600 20.800 125.000 23.100 ;
        RECT 126.200 20.800 126.600 23.100 ;
        RECT 127.800 20.800 128.200 25.100 ;
        RECT 130.600 20.800 131.000 23.100 ;
        RECT 132.200 20.800 132.600 23.100 ;
        RECT 135.000 20.800 135.400 25.000 ;
        RECT 136.900 20.800 137.300 23.100 ;
        RECT 139.000 20.800 139.400 25.100 ;
        RECT 141.400 20.800 141.800 23.100 ;
        RECT 143.000 20.800 143.400 23.100 ;
        RECT 143.800 20.800 144.200 23.100 ;
        RECT 146.200 20.800 146.600 25.100 ;
        RECT 149.000 20.800 149.400 23.100 ;
        RECT 150.600 20.800 151.000 23.100 ;
        RECT 153.400 20.800 153.800 25.000 ;
        RECT 155.000 20.800 155.400 23.100 ;
        RECT 156.600 20.800 157.000 23.100 ;
        RECT 158.200 20.800 158.600 23.100 ;
        RECT 159.800 20.800 160.200 23.100 ;
        RECT 161.400 20.800 161.800 25.000 ;
        RECT 164.200 20.800 164.600 23.100 ;
        RECT 165.800 20.800 166.200 23.100 ;
        RECT 168.600 20.800 169.000 25.100 ;
        RECT 171.000 20.800 171.400 23.100 ;
        RECT 172.100 20.800 172.500 23.100 ;
        RECT 174.200 20.800 174.600 25.100 ;
        RECT 175.000 20.800 175.400 25.100 ;
        RECT 177.100 20.800 177.500 23.100 ;
        RECT 178.200 20.800 178.600 23.100 ;
        RECT 179.800 20.800 180.200 23.100 ;
        RECT 0.200 20.200 180.600 20.800 ;
        RECT 1.200 15.900 1.600 20.200 ;
        RECT 3.800 16.100 4.200 20.200 ;
        RECT 6.200 17.900 6.600 20.200 ;
        RECT 7.800 16.500 8.200 20.200 ;
        RECT 11.800 15.900 12.200 20.200 ;
        RECT 13.400 15.900 13.800 20.200 ;
        RECT 16.200 17.900 16.600 20.200 ;
        RECT 17.800 17.900 18.200 20.200 ;
        RECT 20.600 16.000 21.000 20.200 ;
        RECT 23.000 16.100 23.400 20.200 ;
        RECT 25.600 15.900 26.000 20.200 ;
        RECT 27.800 17.900 28.200 20.200 ;
        RECT 29.400 16.000 29.800 20.200 ;
        RECT 32.200 17.900 32.600 20.200 ;
        RECT 33.800 17.900 34.200 20.200 ;
        RECT 36.600 15.900 37.000 20.200 ;
        RECT 40.600 16.100 41.000 20.200 ;
        RECT 43.200 15.900 43.600 20.200 ;
        RECT 44.600 17.900 45.000 20.200 ;
        RECT 47.000 15.900 47.400 20.200 ;
        RECT 49.800 17.900 50.200 20.200 ;
        RECT 51.400 17.900 51.800 20.200 ;
        RECT 54.200 16.000 54.600 20.200 ;
        RECT 55.800 15.900 56.200 20.200 ;
        RECT 59.800 16.500 60.200 20.200 ;
        RECT 61.400 17.900 61.800 20.200 ;
        RECT 63.600 15.900 64.000 20.200 ;
        RECT 66.200 16.100 66.600 20.200 ;
        RECT 67.800 17.900 68.200 20.200 ;
        RECT 69.400 17.900 69.800 20.200 ;
        RECT 70.200 15.900 70.600 20.200 ;
        RECT 74.200 16.500 74.600 20.200 ;
        RECT 75.800 15.900 76.200 20.200 ;
        RECT 77.400 15.900 77.800 20.200 ;
        RECT 79.000 15.900 79.400 20.200 ;
        RECT 80.600 15.900 81.000 20.200 ;
        RECT 83.400 17.900 83.800 20.200 ;
        RECT 85.000 17.900 85.400 20.200 ;
        RECT 87.800 16.000 88.200 20.200 ;
        RECT 91.000 17.900 91.400 20.200 ;
        RECT 93.200 15.900 93.600 20.200 ;
        RECT 95.800 16.100 96.200 20.200 ;
        RECT 98.200 15.900 98.600 20.200 ;
        RECT 101.000 17.900 101.400 20.200 ;
        RECT 102.600 17.900 103.000 20.200 ;
        RECT 105.400 16.000 105.800 20.200 ;
        RECT 107.000 17.900 107.400 20.200 ;
        RECT 109.200 15.900 109.600 20.200 ;
        RECT 111.800 16.100 112.200 20.200 ;
        RECT 113.400 17.900 113.800 20.200 ;
        RECT 115.800 16.100 116.200 20.200 ;
        RECT 118.400 15.900 118.800 20.200 ;
        RECT 119.800 17.900 120.200 20.200 ;
        RECT 122.200 16.100 122.600 20.200 ;
        RECT 124.800 15.900 125.200 20.200 ;
        RECT 127.000 16.000 127.400 20.200 ;
        RECT 129.800 17.900 130.200 20.200 ;
        RECT 131.400 17.900 131.800 20.200 ;
        RECT 134.200 15.900 134.600 20.200 ;
        RECT 135.800 17.900 136.200 20.200 ;
        RECT 138.000 15.900 138.400 20.200 ;
        RECT 140.600 16.100 141.000 20.200 ;
        RECT 144.400 15.900 144.800 20.200 ;
        RECT 147.000 16.100 147.400 20.200 ;
        RECT 149.400 16.100 149.800 20.200 ;
        RECT 152.000 15.900 152.400 20.200 ;
        RECT 154.200 16.000 154.600 20.200 ;
        RECT 157.000 17.900 157.400 20.200 ;
        RECT 158.600 17.900 159.000 20.200 ;
        RECT 161.400 15.900 161.800 20.200 ;
        RECT 163.800 16.100 164.200 20.200 ;
        RECT 166.400 15.900 166.800 20.200 ;
        RECT 167.800 17.900 168.200 20.200 ;
        RECT 169.400 17.900 169.800 20.200 ;
        RECT 171.000 17.900 171.400 20.200 ;
        RECT 171.800 17.900 172.200 20.200 ;
        RECT 174.200 17.900 174.600 20.200 ;
        RECT 175.600 15.900 176.000 20.200 ;
        RECT 178.200 16.100 178.600 20.200 ;
        RECT 1.400 0.800 1.800 5.000 ;
        RECT 4.200 0.800 4.600 3.100 ;
        RECT 5.800 0.800 6.200 3.100 ;
        RECT 8.600 0.800 9.000 5.100 ;
        RECT 11.000 0.800 11.400 5.000 ;
        RECT 13.800 0.800 14.200 3.100 ;
        RECT 15.400 0.800 15.800 3.100 ;
        RECT 18.200 0.800 18.600 5.100 ;
        RECT 20.600 0.800 21.000 4.500 ;
        RECT 23.000 0.800 23.400 5.100 ;
        RECT 26.200 0.800 26.600 5.000 ;
        RECT 29.000 0.800 29.400 3.100 ;
        RECT 30.600 0.800 31.000 3.100 ;
        RECT 33.400 0.800 33.800 5.100 ;
        RECT 37.400 0.800 37.800 5.000 ;
        RECT 40.200 0.800 40.600 3.100 ;
        RECT 41.800 0.800 42.200 3.100 ;
        RECT 44.600 0.800 45.000 5.100 ;
        RECT 46.200 0.800 46.600 5.100 ;
        RECT 50.200 0.800 50.600 4.500 ;
        RECT 52.600 0.800 53.000 5.000 ;
        RECT 55.400 0.800 55.800 3.100 ;
        RECT 57.000 0.800 57.400 3.100 ;
        RECT 59.800 0.800 60.200 5.100 ;
        RECT 61.400 0.800 61.800 5.100 ;
        RECT 63.000 0.800 63.400 5.100 ;
        RECT 64.600 0.800 65.000 5.100 ;
        RECT 66.200 0.800 66.600 5.100 ;
        RECT 69.000 0.800 69.400 3.100 ;
        RECT 70.600 0.800 71.000 3.100 ;
        RECT 73.400 0.800 73.800 5.000 ;
        RECT 75.800 0.800 76.200 5.000 ;
        RECT 78.600 0.800 79.000 3.100 ;
        RECT 80.200 0.800 80.600 3.100 ;
        RECT 83.000 0.800 83.400 5.100 ;
        RECT 84.600 0.800 85.000 3.100 ;
        RECT 86.800 0.800 87.200 5.100 ;
        RECT 89.400 0.800 89.800 4.900 ;
        RECT 92.600 0.800 93.000 5.100 ;
        RECT 94.200 0.800 94.600 5.100 ;
        RECT 95.800 0.800 96.200 5.100 ;
        RECT 97.400 0.800 97.800 5.100 ;
        RECT 100.200 0.800 100.600 3.100 ;
        RECT 101.800 0.800 102.200 3.100 ;
        RECT 104.600 0.800 105.000 5.000 ;
        RECT 106.200 0.800 106.600 3.100 ;
        RECT 107.800 0.800 108.200 3.100 ;
        RECT 109.400 0.800 109.800 5.000 ;
        RECT 112.200 0.800 112.600 3.100 ;
        RECT 113.800 0.800 114.200 3.100 ;
        RECT 116.600 0.800 117.000 5.100 ;
        RECT 118.200 0.800 118.600 5.100 ;
        RECT 119.800 0.800 120.200 5.100 ;
        RECT 121.400 0.800 121.800 5.100 ;
        RECT 122.200 0.800 122.600 5.100 ;
        RECT 125.400 0.800 125.800 3.100 ;
        RECT 127.000 0.800 127.400 5.000 ;
        RECT 129.800 0.800 130.200 3.100 ;
        RECT 131.400 0.800 131.800 3.100 ;
        RECT 134.200 0.800 134.600 5.100 ;
        RECT 135.800 0.800 136.200 3.100 ;
        RECT 137.400 0.800 137.800 3.100 ;
        RECT 138.200 0.800 138.600 3.100 ;
        RECT 142.000 0.800 142.400 5.100 ;
        RECT 144.600 0.800 145.000 4.900 ;
        RECT 147.000 0.800 147.400 4.900 ;
        RECT 149.600 0.800 150.000 5.100 ;
        RECT 151.800 0.800 152.200 5.000 ;
        RECT 154.600 0.800 155.000 3.100 ;
        RECT 156.200 0.800 156.600 3.100 ;
        RECT 159.000 0.800 159.400 5.100 ;
        RECT 161.400 0.800 161.800 5.000 ;
        RECT 164.200 0.800 164.600 3.100 ;
        RECT 165.800 0.800 166.200 3.100 ;
        RECT 168.600 0.800 169.000 5.100 ;
        RECT 171.000 0.800 171.400 5.000 ;
        RECT 173.800 0.800 174.200 3.100 ;
        RECT 175.400 0.800 175.800 3.100 ;
        RECT 178.200 0.800 178.600 5.100 ;
        RECT 0.200 0.200 180.600 0.800 ;
      LAYER via1 ;
        RECT 131.800 161.800 132.200 162.200 ;
        RECT 139.000 162.700 139.400 163.100 ;
        RECT 37.000 160.300 37.400 160.700 ;
        RECT 37.700 160.300 38.100 160.700 ;
        RECT 138.600 160.300 139.000 160.700 ;
        RECT 139.300 160.300 139.700 160.700 ;
        RECT 159.000 155.600 159.400 156.000 ;
        RECT 165.400 141.800 165.800 142.200 ;
        RECT 37.000 140.300 37.400 140.700 ;
        RECT 37.700 140.300 38.100 140.700 ;
        RECT 138.600 140.300 139.000 140.700 ;
        RECT 139.300 140.300 139.700 140.700 ;
        RECT 37.000 120.300 37.400 120.700 ;
        RECT 37.700 120.300 38.100 120.700 ;
        RECT 138.600 120.300 139.000 120.700 ;
        RECT 139.300 120.300 139.700 120.700 ;
        RECT 37.000 100.300 37.400 100.700 ;
        RECT 37.700 100.300 38.100 100.700 ;
        RECT 138.600 100.300 139.000 100.700 ;
        RECT 139.300 100.300 139.700 100.700 ;
        RECT 138.200 98.800 138.600 99.200 ;
        RECT 131.000 95.600 131.400 96.000 ;
        RECT 138.200 95.800 138.600 96.200 ;
        RECT 144.600 81.800 145.000 82.200 ;
        RECT 37.000 80.300 37.400 80.700 ;
        RECT 37.700 80.300 38.100 80.700 ;
        RECT 138.600 80.300 139.000 80.700 ;
        RECT 139.300 80.300 139.700 80.700 ;
        RECT 151.000 75.600 151.400 76.000 ;
        RECT 37.000 60.300 37.400 60.700 ;
        RECT 37.700 60.300 38.100 60.700 ;
        RECT 138.600 60.300 139.000 60.700 ;
        RECT 139.300 60.300 139.700 60.700 ;
        RECT 37.000 40.300 37.400 40.700 ;
        RECT 37.700 40.300 38.100 40.700 ;
        RECT 138.600 40.300 139.000 40.700 ;
        RECT 139.300 40.300 139.700 40.700 ;
        RECT 37.000 20.300 37.400 20.700 ;
        RECT 37.700 20.300 38.100 20.700 ;
        RECT 138.600 20.300 139.000 20.700 ;
        RECT 139.300 20.300 139.700 20.700 ;
        RECT 37.000 0.300 37.400 0.700 ;
        RECT 37.700 0.300 38.100 0.700 ;
        RECT 138.600 0.300 139.000 0.700 ;
        RECT 139.300 0.300 139.700 0.700 ;
      LAYER metal2 ;
        RECT 131.800 164.800 132.200 165.200 ;
        RECT 139.000 165.000 139.400 165.400 ;
        RECT 131.800 162.200 132.100 164.800 ;
        RECT 139.000 163.100 139.300 165.000 ;
        RECT 139.000 162.700 139.400 163.100 ;
        RECT 131.800 161.800 132.200 162.200 ;
        RECT 36.800 160.300 38.400 160.700 ;
        RECT 138.400 160.300 140.000 160.700 ;
        RECT 159.000 157.900 159.400 158.300 ;
        RECT 159.000 156.000 159.300 157.900 ;
        RECT 159.000 155.600 159.400 156.000 ;
        RECT 165.400 145.000 165.800 145.400 ;
        RECT 165.400 142.200 165.700 145.000 ;
        RECT 165.400 141.800 165.800 142.200 ;
        RECT 36.800 140.300 38.400 140.700 ;
        RECT 138.400 140.300 140.000 140.700 ;
        RECT 36.800 120.300 38.400 120.700 ;
        RECT 138.400 120.300 140.000 120.700 ;
        RECT 36.800 100.300 38.400 100.700 ;
        RECT 138.400 100.300 140.000 100.700 ;
        RECT 138.200 98.800 138.600 99.200 ;
        RECT 131.000 97.900 131.400 98.300 ;
        RECT 131.000 96.000 131.300 97.900 ;
        RECT 138.200 96.200 138.500 98.800 ;
        RECT 131.000 95.600 131.400 96.000 ;
        RECT 138.200 95.800 138.600 96.200 ;
        RECT 144.600 85.000 145.000 85.400 ;
        RECT 144.600 82.200 144.900 85.000 ;
        RECT 144.600 81.800 145.000 82.200 ;
        RECT 36.800 80.300 38.400 80.700 ;
        RECT 138.400 80.300 140.000 80.700 ;
        RECT 151.000 77.900 151.400 78.300 ;
        RECT 151.000 76.000 151.300 77.900 ;
        RECT 151.000 75.600 151.400 76.000 ;
        RECT 36.800 60.300 38.400 60.700 ;
        RECT 138.400 60.300 140.000 60.700 ;
        RECT 36.800 40.300 38.400 40.700 ;
        RECT 138.400 40.300 140.000 40.700 ;
        RECT 36.800 20.300 38.400 20.700 ;
        RECT 138.400 20.300 140.000 20.700 ;
        RECT 36.800 0.300 38.400 0.700 ;
        RECT 138.400 0.300 140.000 0.700 ;
      LAYER via2 ;
        RECT 37.000 160.300 37.400 160.700 ;
        RECT 37.700 160.300 38.100 160.700 ;
        RECT 138.600 160.300 139.000 160.700 ;
        RECT 139.300 160.300 139.700 160.700 ;
        RECT 37.000 140.300 37.400 140.700 ;
        RECT 37.700 140.300 38.100 140.700 ;
        RECT 138.600 140.300 139.000 140.700 ;
        RECT 139.300 140.300 139.700 140.700 ;
        RECT 37.000 120.300 37.400 120.700 ;
        RECT 37.700 120.300 38.100 120.700 ;
        RECT 138.600 120.300 139.000 120.700 ;
        RECT 139.300 120.300 139.700 120.700 ;
        RECT 37.000 100.300 37.400 100.700 ;
        RECT 37.700 100.300 38.100 100.700 ;
        RECT 138.600 100.300 139.000 100.700 ;
        RECT 139.300 100.300 139.700 100.700 ;
        RECT 37.000 80.300 37.400 80.700 ;
        RECT 37.700 80.300 38.100 80.700 ;
        RECT 138.600 80.300 139.000 80.700 ;
        RECT 139.300 80.300 139.700 80.700 ;
        RECT 37.000 60.300 37.400 60.700 ;
        RECT 37.700 60.300 38.100 60.700 ;
        RECT 138.600 60.300 139.000 60.700 ;
        RECT 139.300 60.300 139.700 60.700 ;
        RECT 37.000 40.300 37.400 40.700 ;
        RECT 37.700 40.300 38.100 40.700 ;
        RECT 138.600 40.300 139.000 40.700 ;
        RECT 139.300 40.300 139.700 40.700 ;
        RECT 37.000 20.300 37.400 20.700 ;
        RECT 37.700 20.300 38.100 20.700 ;
        RECT 138.600 20.300 139.000 20.700 ;
        RECT 139.300 20.300 139.700 20.700 ;
        RECT 37.000 0.300 37.400 0.700 ;
        RECT 37.700 0.300 38.100 0.700 ;
        RECT 138.600 0.300 139.000 0.700 ;
        RECT 139.300 0.300 139.700 0.700 ;
      LAYER metal3 ;
        RECT 36.800 160.300 38.400 160.700 ;
        RECT 138.400 160.300 140.000 160.700 ;
        RECT 36.800 140.300 38.400 140.700 ;
        RECT 138.400 140.300 140.000 140.700 ;
        RECT 36.800 120.300 38.400 120.700 ;
        RECT 138.400 120.300 140.000 120.700 ;
        RECT 36.800 100.300 38.400 100.700 ;
        RECT 138.400 100.300 140.000 100.700 ;
        RECT 36.800 80.300 38.400 80.700 ;
        RECT 138.400 80.300 140.000 80.700 ;
        RECT 36.800 60.300 38.400 60.700 ;
        RECT 138.400 60.300 140.000 60.700 ;
        RECT 36.800 40.300 38.400 40.700 ;
        RECT 138.400 40.300 140.000 40.700 ;
        RECT 36.800 20.300 38.400 20.700 ;
        RECT 138.400 20.300 140.000 20.700 ;
        RECT 36.800 0.300 38.400 0.700 ;
        RECT 138.400 0.300 140.000 0.700 ;
      LAYER via3 ;
        RECT 37.000 160.300 37.400 160.700 ;
        RECT 37.800 160.300 38.200 160.700 ;
        RECT 138.600 160.300 139.000 160.700 ;
        RECT 139.400 160.300 139.800 160.700 ;
        RECT 37.000 140.300 37.400 140.700 ;
        RECT 37.800 140.300 38.200 140.700 ;
        RECT 138.600 140.300 139.000 140.700 ;
        RECT 139.400 140.300 139.800 140.700 ;
        RECT 37.000 120.300 37.400 120.700 ;
        RECT 37.800 120.300 38.200 120.700 ;
        RECT 138.600 120.300 139.000 120.700 ;
        RECT 139.400 120.300 139.800 120.700 ;
        RECT 37.000 100.300 37.400 100.700 ;
        RECT 37.800 100.300 38.200 100.700 ;
        RECT 138.600 100.300 139.000 100.700 ;
        RECT 139.400 100.300 139.800 100.700 ;
        RECT 37.000 80.300 37.400 80.700 ;
        RECT 37.800 80.300 38.200 80.700 ;
        RECT 138.600 80.300 139.000 80.700 ;
        RECT 139.400 80.300 139.800 80.700 ;
        RECT 37.000 60.300 37.400 60.700 ;
        RECT 37.800 60.300 38.200 60.700 ;
        RECT 138.600 60.300 139.000 60.700 ;
        RECT 139.400 60.300 139.800 60.700 ;
        RECT 37.000 40.300 37.400 40.700 ;
        RECT 37.800 40.300 38.200 40.700 ;
        RECT 138.600 40.300 139.000 40.700 ;
        RECT 139.400 40.300 139.800 40.700 ;
        RECT 37.000 20.300 37.400 20.700 ;
        RECT 37.800 20.300 38.200 20.700 ;
        RECT 138.600 20.300 139.000 20.700 ;
        RECT 139.400 20.300 139.800 20.700 ;
        RECT 37.000 0.300 37.400 0.700 ;
        RECT 37.800 0.300 38.200 0.700 ;
        RECT 138.600 0.300 139.000 0.700 ;
        RECT 139.400 0.300 139.800 0.700 ;
      LAYER metal4 ;
        RECT 36.800 160.300 38.400 160.700 ;
        RECT 138.400 160.300 140.000 160.700 ;
        RECT 36.800 140.300 38.400 140.700 ;
        RECT 138.400 140.300 140.000 140.700 ;
        RECT 36.800 120.300 38.400 120.700 ;
        RECT 138.400 120.300 140.000 120.700 ;
        RECT 36.800 100.300 38.400 100.700 ;
        RECT 138.400 100.300 140.000 100.700 ;
        RECT 36.800 80.300 38.400 80.700 ;
        RECT 138.400 80.300 140.000 80.700 ;
        RECT 36.800 60.300 38.400 60.700 ;
        RECT 138.400 60.300 140.000 60.700 ;
        RECT 36.800 40.300 38.400 40.700 ;
        RECT 138.400 40.300 140.000 40.700 ;
        RECT 36.800 20.300 38.400 20.700 ;
        RECT 138.400 20.300 140.000 20.700 ;
        RECT 36.800 0.300 38.400 0.700 ;
        RECT 138.400 0.300 140.000 0.700 ;
      LAYER via4 ;
        RECT 37.000 160.300 37.400 160.700 ;
        RECT 37.700 160.300 38.100 160.700 ;
        RECT 138.600 160.300 139.000 160.700 ;
        RECT 139.300 160.300 139.700 160.700 ;
        RECT 37.000 140.300 37.400 140.700 ;
        RECT 37.700 140.300 38.100 140.700 ;
        RECT 138.600 140.300 139.000 140.700 ;
        RECT 139.300 140.300 139.700 140.700 ;
        RECT 37.000 120.300 37.400 120.700 ;
        RECT 37.700 120.300 38.100 120.700 ;
        RECT 138.600 120.300 139.000 120.700 ;
        RECT 139.300 120.300 139.700 120.700 ;
        RECT 37.000 100.300 37.400 100.700 ;
        RECT 37.700 100.300 38.100 100.700 ;
        RECT 138.600 100.300 139.000 100.700 ;
        RECT 139.300 100.300 139.700 100.700 ;
        RECT 37.000 80.300 37.400 80.700 ;
        RECT 37.700 80.300 38.100 80.700 ;
        RECT 138.600 80.300 139.000 80.700 ;
        RECT 139.300 80.300 139.700 80.700 ;
        RECT 37.000 60.300 37.400 60.700 ;
        RECT 37.700 60.300 38.100 60.700 ;
        RECT 138.600 60.300 139.000 60.700 ;
        RECT 139.300 60.300 139.700 60.700 ;
        RECT 37.000 40.300 37.400 40.700 ;
        RECT 37.700 40.300 38.100 40.700 ;
        RECT 138.600 40.300 139.000 40.700 ;
        RECT 139.300 40.300 139.700 40.700 ;
        RECT 37.000 20.300 37.400 20.700 ;
        RECT 37.700 20.300 38.100 20.700 ;
        RECT 138.600 20.300 139.000 20.700 ;
        RECT 139.300 20.300 139.700 20.700 ;
        RECT 37.000 0.300 37.400 0.700 ;
        RECT 37.700 0.300 38.100 0.700 ;
        RECT 138.600 0.300 139.000 0.700 ;
        RECT 139.300 0.300 139.700 0.700 ;
      LAYER metal5 ;
        RECT 36.800 160.200 38.400 160.700 ;
        RECT 138.400 160.200 140.000 160.700 ;
        RECT 36.800 140.200 38.400 140.700 ;
        RECT 138.400 140.200 140.000 140.700 ;
        RECT 36.800 120.200 38.400 120.700 ;
        RECT 138.400 120.200 140.000 120.700 ;
        RECT 36.800 100.200 38.400 100.700 ;
        RECT 138.400 100.200 140.000 100.700 ;
        RECT 36.800 80.200 38.400 80.700 ;
        RECT 138.400 80.200 140.000 80.700 ;
        RECT 36.800 60.200 38.400 60.700 ;
        RECT 138.400 60.200 140.000 60.700 ;
        RECT 36.800 40.200 38.400 40.700 ;
        RECT 138.400 40.200 140.000 40.700 ;
        RECT 36.800 20.200 38.400 20.700 ;
        RECT 138.400 20.200 140.000 20.700 ;
        RECT 36.800 0.200 38.400 0.700 ;
        RECT 138.400 0.200 140.000 0.700 ;
      LAYER via5 ;
        RECT 37.800 160.200 38.300 160.700 ;
        RECT 139.400 160.200 139.900 160.700 ;
        RECT 37.800 140.200 38.300 140.700 ;
        RECT 139.400 140.200 139.900 140.700 ;
        RECT 37.800 120.200 38.300 120.700 ;
        RECT 139.400 120.200 139.900 120.700 ;
        RECT 37.800 100.200 38.300 100.700 ;
        RECT 139.400 100.200 139.900 100.700 ;
        RECT 37.800 80.200 38.300 80.700 ;
        RECT 139.400 80.200 139.900 80.700 ;
        RECT 37.800 60.200 38.300 60.700 ;
        RECT 139.400 60.200 139.900 60.700 ;
        RECT 37.800 40.200 38.300 40.700 ;
        RECT 139.400 40.200 139.900 40.700 ;
        RECT 37.800 20.200 38.300 20.700 ;
        RECT 139.400 20.200 139.900 20.700 ;
        RECT 37.800 0.200 38.300 0.700 ;
        RECT 139.400 0.200 139.900 0.700 ;
      LAYER metal6 ;
        RECT 36.800 -3.000 38.400 173.000 ;
        RECT 138.400 -3.000 140.000 173.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 170.200 180.600 170.800 ;
        RECT 1.400 168.900 1.800 170.200 ;
        RECT 2.800 167.500 3.200 170.200 ;
        RECT 5.400 167.700 5.800 170.200 ;
        RECT 7.800 167.900 8.200 170.200 ;
        RECT 10.500 168.900 11.000 170.200 ;
        RECT 12.200 168.900 12.600 170.200 ;
        RECT 15.000 168.000 15.400 170.200 ;
        RECT 17.400 167.900 17.800 170.200 ;
        RECT 20.100 168.900 20.600 170.200 ;
        RECT 21.800 168.900 22.200 170.200 ;
        RECT 24.600 168.000 25.000 170.200 ;
        RECT 27.000 168.000 27.400 170.200 ;
        RECT 29.800 168.900 30.200 170.200 ;
        RECT 31.400 168.900 31.900 170.200 ;
        RECT 34.200 167.900 34.600 170.200 ;
        RECT 38.200 167.700 38.600 170.200 ;
        RECT 40.800 167.500 41.200 170.200 ;
        RECT 43.000 168.900 43.400 170.200 ;
        RECT 44.600 167.900 45.000 170.200 ;
        RECT 47.300 168.900 47.800 170.200 ;
        RECT 49.000 168.900 49.400 170.200 ;
        RECT 51.800 168.000 52.200 170.200 ;
        RECT 53.400 167.900 53.800 170.200 ;
        RECT 55.000 167.900 55.400 170.200 ;
        RECT 56.600 167.900 57.000 170.200 ;
        RECT 58.200 167.900 58.600 170.200 ;
        RECT 59.800 167.900 60.200 170.200 ;
        RECT 61.400 167.900 61.800 170.200 ;
        RECT 64.100 168.900 64.600 170.200 ;
        RECT 65.800 168.900 66.200 170.200 ;
        RECT 68.600 168.000 69.000 170.200 ;
        RECT 70.200 167.900 70.600 170.200 ;
        RECT 71.800 167.900 72.200 170.200 ;
        RECT 73.400 167.900 73.800 170.200 ;
        RECT 74.200 167.900 74.600 170.200 ;
        RECT 75.800 167.900 76.200 170.200 ;
        RECT 77.400 167.900 77.800 170.200 ;
        RECT 79.000 167.900 79.400 170.200 ;
        RECT 80.600 167.900 81.000 170.200 ;
        RECT 81.400 167.900 81.800 170.200 ;
        RECT 83.000 167.900 83.400 170.200 ;
        RECT 84.600 167.900 85.000 170.200 ;
        RECT 85.400 167.900 85.800 170.200 ;
        RECT 87.000 167.900 87.400 170.200 ;
        RECT 88.600 167.900 89.000 170.200 ;
        RECT 91.800 167.900 92.200 170.200 ;
        RECT 94.500 168.900 95.000 170.200 ;
        RECT 96.200 168.900 96.600 170.200 ;
        RECT 99.000 168.000 99.400 170.200 ;
        RECT 101.400 167.700 101.800 170.200 ;
        RECT 104.000 167.500 104.400 170.200 ;
        RECT 106.200 168.900 106.600 170.200 ;
        RECT 107.800 168.000 108.200 170.200 ;
        RECT 110.600 168.900 111.000 170.200 ;
        RECT 112.200 168.900 112.700 170.200 ;
        RECT 115.000 167.900 115.400 170.200 ;
        RECT 116.600 168.900 117.000 170.200 ;
        RECT 119.800 167.900 120.200 170.200 ;
        RECT 125.400 168.900 125.800 170.200 ;
        RECT 127.000 168.900 127.400 170.200 ;
        RECT 131.800 167.900 132.200 170.200 ;
        RECT 137.400 167.900 137.800 170.200 ;
        RECT 142.200 168.900 142.600 170.200 ;
        RECT 143.800 168.900 144.200 170.200 ;
        RECT 149.400 167.900 149.800 170.200 ;
        RECT 152.600 168.900 153.000 170.200 ;
        RECT 154.200 167.900 154.600 170.200 ;
        RECT 156.600 167.900 157.000 170.200 ;
        RECT 159.300 168.900 159.800 170.200 ;
        RECT 161.000 168.900 161.400 170.200 ;
        RECT 163.800 168.000 164.200 170.200 ;
        RECT 166.200 167.700 166.600 170.200 ;
        RECT 168.800 167.500 169.200 170.200 ;
        RECT 171.000 167.700 171.400 170.200 ;
        RECT 173.600 167.500 174.000 170.200 ;
        RECT 175.800 167.900 176.200 170.200 ;
        RECT 178.200 167.900 178.600 170.200 ;
        RECT 1.400 150.800 1.800 153.100 ;
        RECT 4.100 150.800 4.600 152.100 ;
        RECT 5.800 150.800 6.200 152.100 ;
        RECT 8.600 150.800 9.000 153.000 ;
        RECT 10.200 150.800 10.600 152.100 ;
        RECT 12.400 150.800 12.800 153.500 ;
        RECT 15.000 150.800 15.400 153.300 ;
        RECT 16.600 150.800 17.000 153.100 ;
        RECT 19.800 150.800 20.200 153.300 ;
        RECT 22.400 150.800 22.800 153.500 ;
        RECT 24.600 150.800 25.000 152.100 ;
        RECT 25.400 150.800 25.800 153.100 ;
        RECT 27.800 150.800 28.200 153.100 ;
        RECT 29.400 150.800 29.800 153.100 ;
        RECT 31.000 150.800 31.400 153.100 ;
        RECT 32.600 150.800 33.000 153.100 ;
        RECT 34.200 150.800 34.600 153.100 ;
        RECT 37.400 150.800 37.800 153.100 ;
        RECT 40.100 150.800 40.600 152.100 ;
        RECT 41.800 150.800 42.200 152.100 ;
        RECT 44.600 150.800 45.000 153.000 ;
        RECT 46.200 150.800 46.600 152.100 ;
        RECT 47.800 150.800 48.200 152.100 ;
        RECT 48.600 150.800 49.000 152.100 ;
        RECT 50.700 150.800 51.100 153.100 ;
        RECT 52.600 150.800 53.000 153.300 ;
        RECT 55.200 150.800 55.600 153.500 ;
        RECT 57.400 150.800 57.800 152.100 ;
        RECT 58.200 150.800 58.600 153.100 ;
        RECT 61.400 150.800 61.800 153.300 ;
        RECT 64.000 150.800 64.400 153.500 ;
        RECT 66.200 150.800 66.600 152.100 ;
        RECT 67.800 150.800 68.200 153.000 ;
        RECT 70.600 150.800 71.000 152.100 ;
        RECT 72.200 150.800 72.700 152.100 ;
        RECT 75.000 150.800 75.400 153.100 ;
        RECT 76.900 150.800 77.300 153.100 ;
        RECT 79.000 150.800 79.400 152.100 ;
        RECT 80.600 150.800 81.000 153.100 ;
        RECT 83.300 150.800 83.800 152.100 ;
        RECT 85.000 150.800 85.400 152.100 ;
        RECT 87.800 150.800 88.200 153.000 ;
        RECT 91.800 150.800 92.200 153.300 ;
        RECT 94.400 150.800 94.800 153.500 ;
        RECT 96.600 150.800 97.000 152.100 ;
        RECT 97.400 150.800 97.800 152.100 ;
        RECT 99.600 150.800 100.000 153.500 ;
        RECT 102.200 150.800 102.600 153.300 ;
        RECT 104.600 150.800 105.000 153.000 ;
        RECT 107.400 150.800 107.800 152.100 ;
        RECT 109.000 150.800 109.500 152.100 ;
        RECT 111.800 150.800 112.200 153.100 ;
        RECT 114.200 150.800 114.600 153.000 ;
        RECT 117.000 150.800 117.400 152.100 ;
        RECT 118.600 150.800 119.100 152.100 ;
        RECT 121.400 150.800 121.800 153.100 ;
        RECT 123.000 150.800 123.400 152.100 ;
        RECT 125.200 150.800 125.600 153.500 ;
        RECT 127.800 150.800 128.200 153.300 ;
        RECT 130.200 150.800 130.600 153.300 ;
        RECT 132.800 150.800 133.200 153.500 ;
        RECT 135.000 150.800 135.400 152.100 ;
        RECT 138.200 150.800 138.600 153.100 ;
        RECT 140.900 150.800 141.400 152.100 ;
        RECT 142.600 150.800 143.000 152.100 ;
        RECT 145.400 150.800 145.800 153.000 ;
        RECT 147.000 150.800 147.400 153.100 ;
        RECT 148.600 150.800 149.000 153.100 ;
        RECT 150.200 150.800 150.600 153.100 ;
        RECT 151.800 150.800 152.200 153.100 ;
        RECT 153.400 150.800 153.800 153.100 ;
        RECT 154.200 150.800 154.600 152.100 ;
        RECT 157.400 150.800 157.800 153.100 ;
        RECT 162.200 150.800 162.600 152.100 ;
        RECT 163.800 150.800 164.200 152.100 ;
        RECT 169.400 150.800 169.800 153.100 ;
        RECT 172.600 150.800 173.000 152.100 ;
        RECT 174.200 150.800 174.600 153.100 ;
        RECT 176.600 150.800 177.000 152.100 ;
        RECT 178.200 150.800 178.600 153.100 ;
        RECT 0.200 150.200 180.600 150.800 ;
        RECT 1.400 147.900 1.800 150.200 ;
        RECT 4.100 148.900 4.600 150.200 ;
        RECT 5.800 148.900 6.200 150.200 ;
        RECT 8.600 148.000 9.000 150.200 ;
        RECT 10.200 148.900 10.600 150.200 ;
        RECT 11.800 148.900 12.200 150.200 ;
        RECT 12.600 148.900 13.000 150.200 ;
        RECT 14.700 147.900 15.100 150.200 ;
        RECT 15.800 147.900 16.200 150.200 ;
        RECT 18.200 146.900 18.600 150.200 ;
        RECT 22.200 147.700 22.600 150.200 ;
        RECT 24.800 147.500 25.200 150.200 ;
        RECT 27.000 148.900 27.400 150.200 ;
        RECT 28.600 148.000 29.000 150.200 ;
        RECT 31.400 148.900 31.800 150.200 ;
        RECT 33.000 148.900 33.500 150.200 ;
        RECT 35.800 147.900 36.200 150.200 ;
        RECT 39.300 147.900 39.700 150.200 ;
        RECT 41.400 148.900 41.800 150.200 ;
        RECT 42.200 148.900 42.600 150.200 ;
        RECT 43.800 148.900 44.200 150.200 ;
        RECT 44.600 147.900 45.000 150.200 ;
        RECT 47.800 147.900 48.200 150.200 ;
        RECT 50.500 148.900 51.000 150.200 ;
        RECT 52.200 148.900 52.600 150.200 ;
        RECT 55.000 148.000 55.400 150.200 ;
        RECT 59.000 146.900 59.400 150.200 ;
        RECT 59.800 147.900 60.200 150.200 ;
        RECT 63.000 148.900 63.400 150.200 ;
        RECT 64.600 149.100 65.000 150.200 ;
        RECT 69.400 148.000 69.800 150.200 ;
        RECT 72.200 148.900 72.600 150.200 ;
        RECT 73.800 148.900 74.300 150.200 ;
        RECT 76.600 147.900 77.000 150.200 ;
        RECT 78.200 148.900 78.600 150.200 ;
        RECT 79.800 148.900 80.200 150.200 ;
        RECT 81.400 147.700 81.800 150.200 ;
        RECT 84.000 147.500 84.400 150.200 ;
        RECT 86.200 148.900 86.600 150.200 ;
        RECT 89.400 148.000 89.800 150.200 ;
        RECT 92.200 148.900 92.600 150.200 ;
        RECT 93.800 148.900 94.300 150.200 ;
        RECT 96.600 147.900 97.000 150.200 ;
        RECT 99.800 147.900 100.200 150.200 ;
        RECT 100.600 147.900 101.000 150.200 ;
        RECT 103.600 147.900 104.000 150.200 ;
        RECT 104.800 147.900 105.200 150.200 ;
        RECT 107.800 147.900 108.200 150.200 ;
        RECT 108.600 148.900 109.000 150.200 ;
        RECT 110.800 147.500 111.200 150.200 ;
        RECT 113.400 147.700 113.800 150.200 ;
        RECT 115.800 147.700 116.200 150.200 ;
        RECT 118.400 147.500 118.800 150.200 ;
        RECT 120.600 148.900 121.000 150.200 ;
        RECT 122.200 148.000 122.600 150.200 ;
        RECT 125.000 148.900 125.400 150.200 ;
        RECT 126.600 148.900 127.100 150.200 ;
        RECT 129.400 147.900 129.800 150.200 ;
        RECT 131.600 147.500 132.000 150.200 ;
        RECT 134.200 147.700 134.600 150.200 ;
        RECT 136.600 148.900 137.000 150.200 ;
        RECT 139.800 148.000 140.200 150.200 ;
        RECT 142.600 148.900 143.000 150.200 ;
        RECT 144.200 148.900 144.700 150.200 ;
        RECT 147.000 147.900 147.400 150.200 ;
        RECT 148.900 147.900 149.300 150.200 ;
        RECT 151.000 148.900 151.400 150.200 ;
        RECT 151.800 148.900 152.200 150.200 ;
        RECT 153.400 148.900 153.800 150.200 ;
        RECT 154.200 148.900 154.600 150.200 ;
        RECT 155.800 148.900 156.200 150.200 ;
        RECT 156.900 147.900 157.300 150.200 ;
        RECT 159.000 148.900 159.400 150.200 ;
        RECT 159.800 148.900 160.200 150.200 ;
        RECT 161.400 148.900 161.800 150.200 ;
        RECT 163.800 147.900 164.200 150.200 ;
        RECT 168.600 148.900 169.000 150.200 ;
        RECT 170.200 148.900 170.600 150.200 ;
        RECT 175.800 147.900 176.200 150.200 ;
        RECT 179.000 148.900 179.400 150.200 ;
        RECT 1.400 130.800 1.800 133.100 ;
        RECT 4.100 130.800 4.600 132.100 ;
        RECT 5.800 130.800 6.200 132.100 ;
        RECT 8.600 130.800 9.000 133.000 ;
        RECT 11.000 130.800 11.400 133.100 ;
        RECT 13.700 130.800 14.200 132.100 ;
        RECT 15.400 130.800 15.800 132.100 ;
        RECT 18.200 130.800 18.600 133.000 ;
        RECT 20.600 130.800 21.000 133.300 ;
        RECT 23.200 130.800 23.600 133.500 ;
        RECT 25.400 130.800 25.800 132.100 ;
        RECT 26.200 130.800 26.600 134.100 ;
        RECT 29.400 130.800 29.800 133.100 ;
        RECT 31.800 130.800 32.200 134.100 ;
        RECT 35.000 130.800 35.400 134.100 ;
        RECT 40.600 130.800 41.000 133.100 ;
        RECT 43.300 130.800 43.800 132.100 ;
        RECT 45.000 130.800 45.400 132.100 ;
        RECT 47.800 130.800 48.200 133.000 ;
        RECT 49.400 130.800 49.800 132.100 ;
        RECT 51.000 130.800 51.400 132.100 ;
        RECT 51.800 130.800 52.200 132.100 ;
        RECT 53.900 130.800 54.300 133.100 ;
        RECT 55.000 130.800 55.400 134.100 ;
        RECT 58.200 130.800 58.600 133.100 ;
        RECT 60.600 130.800 61.000 134.100 ;
        RECT 63.800 130.800 64.200 133.100 ;
        RECT 67.800 130.800 68.200 133.100 ;
        RECT 68.600 130.800 69.000 133.100 ;
        RECT 71.800 130.800 72.200 132.100 ;
        RECT 73.400 130.800 73.800 133.300 ;
        RECT 76.000 130.800 76.400 133.500 ;
        RECT 79.000 130.800 79.400 133.100 ;
        RECT 81.400 130.800 81.800 133.100 ;
        RECT 83.000 130.800 83.400 132.100 ;
        RECT 84.600 130.800 85.000 131.900 ;
        RECT 90.200 130.800 90.600 133.100 ;
        RECT 92.800 130.800 93.200 133.100 ;
        RECT 95.800 130.800 96.200 133.100 ;
        RECT 97.400 130.800 97.800 133.000 ;
        RECT 100.200 130.800 100.600 132.100 ;
        RECT 101.800 130.800 102.300 132.100 ;
        RECT 104.600 130.800 105.000 133.100 ;
        RECT 106.400 130.800 106.800 133.100 ;
        RECT 109.400 130.800 109.800 133.100 ;
        RECT 110.200 130.800 110.600 132.100 ;
        RECT 112.400 130.800 112.800 133.500 ;
        RECT 115.000 130.800 115.400 133.300 ;
        RECT 117.400 130.800 117.800 133.100 ;
        RECT 120.100 130.800 120.600 132.100 ;
        RECT 121.800 130.800 122.200 132.100 ;
        RECT 124.600 130.800 125.000 133.000 ;
        RECT 126.200 130.800 126.600 132.100 ;
        RECT 128.400 130.800 128.800 133.500 ;
        RECT 131.000 130.800 131.400 133.300 ;
        RECT 133.200 130.800 133.600 133.500 ;
        RECT 135.800 130.800 136.200 133.300 ;
        RECT 139.800 130.800 140.200 133.000 ;
        RECT 142.600 130.800 143.000 132.100 ;
        RECT 144.200 130.800 144.700 132.100 ;
        RECT 147.000 130.800 147.400 133.100 ;
        RECT 150.200 130.800 150.600 132.700 ;
        RECT 151.800 130.800 152.200 132.100 ;
        RECT 154.000 130.800 154.400 133.500 ;
        RECT 156.600 130.800 157.000 133.300 ;
        RECT 159.000 130.800 159.400 132.100 ;
        RECT 160.600 130.800 161.000 131.900 ;
        RECT 166.200 130.800 166.600 132.700 ;
        RECT 168.600 130.800 169.000 133.300 ;
        RECT 171.200 130.800 171.600 133.500 ;
        RECT 173.400 130.800 173.800 133.300 ;
        RECT 176.000 130.800 176.400 133.500 ;
        RECT 178.200 130.800 178.600 132.100 ;
        RECT 179.800 130.800 180.200 132.100 ;
        RECT 0.200 130.200 180.600 130.800 ;
        RECT 1.200 127.500 1.600 130.200 ;
        RECT 3.800 127.700 4.200 130.200 ;
        RECT 6.200 128.900 6.600 130.200 ;
        RECT 7.800 127.700 8.200 130.200 ;
        RECT 10.400 127.500 10.800 130.200 ;
        RECT 12.600 128.900 13.000 130.200 ;
        RECT 14.200 127.900 14.600 130.200 ;
        RECT 16.900 128.900 17.400 130.200 ;
        RECT 18.600 128.900 19.000 130.200 ;
        RECT 21.400 128.000 21.800 130.200 ;
        RECT 23.000 126.900 23.400 130.200 ;
        RECT 27.000 127.900 27.400 130.200 ;
        RECT 29.700 128.900 30.200 130.200 ;
        RECT 31.400 128.900 31.800 130.200 ;
        RECT 34.200 128.000 34.600 130.200 ;
        RECT 38.200 127.700 38.600 130.200 ;
        RECT 40.800 127.500 41.200 130.200 ;
        RECT 43.000 128.900 43.400 130.200 ;
        RECT 44.600 127.700 45.000 130.200 ;
        RECT 47.200 127.500 47.600 130.200 ;
        RECT 49.400 128.900 49.800 130.200 ;
        RECT 51.000 127.900 51.400 130.200 ;
        RECT 53.700 128.900 54.200 130.200 ;
        RECT 55.400 128.900 55.800 130.200 ;
        RECT 58.200 128.000 58.600 130.200 ;
        RECT 62.200 126.900 62.600 130.200 ;
        RECT 63.000 126.900 63.400 130.200 ;
        RECT 68.600 126.900 69.000 130.200 ;
        RECT 69.400 126.900 69.800 130.200 ;
        RECT 72.600 126.900 73.000 130.200 ;
        RECT 76.600 128.900 77.000 130.200 ;
        RECT 78.200 129.100 78.600 130.200 ;
        RECT 83.000 127.900 83.400 130.200 ;
        RECT 85.700 128.900 86.200 130.200 ;
        RECT 87.400 128.900 87.800 130.200 ;
        RECT 90.200 128.000 90.600 130.200 ;
        RECT 93.400 128.900 93.800 130.200 ;
        RECT 95.600 127.500 96.000 130.200 ;
        RECT 98.200 127.700 98.600 130.200 ;
        RECT 101.400 127.900 101.800 130.200 ;
        RECT 102.500 127.900 102.900 130.200 ;
        RECT 104.600 128.900 105.000 130.200 ;
        RECT 105.400 128.900 105.800 130.200 ;
        RECT 107.000 128.900 107.400 130.200 ;
        RECT 108.600 128.000 109.000 130.200 ;
        RECT 111.400 128.900 111.800 130.200 ;
        RECT 113.000 128.900 113.500 130.200 ;
        RECT 115.800 127.900 116.200 130.200 ;
        RECT 118.200 128.000 118.600 130.200 ;
        RECT 121.000 128.900 121.400 130.200 ;
        RECT 122.600 128.900 123.100 130.200 ;
        RECT 125.400 127.900 125.800 130.200 ;
        RECT 127.000 128.900 127.400 130.200 ;
        RECT 129.400 127.700 129.800 130.200 ;
        RECT 132.000 127.500 132.400 130.200 ;
        RECT 135.800 128.300 136.200 130.200 ;
        RECT 138.200 128.900 138.600 130.200 ;
        RECT 140.900 127.900 141.300 130.200 ;
        RECT 143.000 128.900 143.400 130.200 ;
        RECT 147.000 129.100 147.400 130.200 ;
        RECT 148.600 128.900 149.000 130.200 ;
        RECT 151.000 128.000 151.400 130.200 ;
        RECT 153.800 128.900 154.200 130.200 ;
        RECT 155.400 128.900 155.900 130.200 ;
        RECT 158.200 127.900 158.600 130.200 ;
        RECT 162.200 128.300 162.600 130.200 ;
        RECT 164.600 127.700 165.000 130.200 ;
        RECT 167.200 127.500 167.600 130.200 ;
        RECT 168.600 128.900 169.000 130.200 ;
        RECT 170.200 128.900 170.600 130.200 ;
        RECT 171.800 127.900 172.200 130.200 ;
        RECT 174.500 128.900 175.000 130.200 ;
        RECT 176.200 128.900 176.600 130.200 ;
        RECT 179.000 128.000 179.400 130.200 ;
        RECT 1.200 110.800 1.600 113.500 ;
        RECT 3.800 110.800 4.200 113.300 ;
        RECT 6.200 110.800 6.600 112.100 ;
        RECT 7.800 110.800 8.200 113.100 ;
        RECT 10.500 110.800 11.000 112.100 ;
        RECT 12.200 110.800 12.600 112.100 ;
        RECT 15.000 110.800 15.400 113.000 ;
        RECT 16.900 110.800 17.300 113.100 ;
        RECT 19.000 110.800 19.400 112.100 ;
        RECT 19.800 110.800 20.200 112.100 ;
        RECT 21.400 110.800 21.800 112.100 ;
        RECT 23.000 110.800 23.400 113.100 ;
        RECT 25.700 110.800 26.200 112.100 ;
        RECT 27.400 110.800 27.800 112.100 ;
        RECT 30.200 110.800 30.600 113.000 ;
        RECT 32.100 110.800 32.500 113.100 ;
        RECT 34.200 110.800 34.600 112.100 ;
        RECT 35.000 110.800 35.400 112.100 ;
        RECT 36.600 110.800 37.000 112.100 ;
        RECT 39.000 110.800 39.400 113.100 ;
        RECT 42.200 110.800 42.600 113.300 ;
        RECT 44.800 110.800 45.200 113.500 ;
        RECT 47.000 110.800 47.400 112.100 ;
        RECT 48.600 110.800 49.000 113.100 ;
        RECT 51.300 110.800 51.800 112.100 ;
        RECT 53.000 110.800 53.400 112.100 ;
        RECT 55.800 110.800 56.200 113.000 ;
        RECT 58.200 110.800 58.600 113.000 ;
        RECT 61.000 110.800 61.400 112.100 ;
        RECT 62.600 110.800 63.100 112.100 ;
        RECT 65.400 110.800 65.800 113.100 ;
        RECT 67.000 110.800 67.400 112.100 ;
        RECT 69.200 110.800 69.600 113.500 ;
        RECT 71.800 110.800 72.200 113.300 ;
        RECT 74.200 110.800 74.600 112.100 ;
        RECT 75.800 110.800 76.200 111.900 ;
        RECT 82.200 110.800 82.600 114.100 ;
        RECT 84.600 110.800 85.000 113.100 ;
        RECT 86.200 110.800 86.600 113.300 ;
        RECT 88.800 110.800 89.200 113.500 ;
        RECT 92.600 110.800 93.000 112.100 ;
        RECT 93.600 110.800 94.000 113.100 ;
        RECT 96.600 110.800 97.000 113.100 ;
        RECT 99.000 110.800 99.400 113.100 ;
        RECT 100.600 110.800 101.000 113.000 ;
        RECT 103.400 110.800 103.800 112.100 ;
        RECT 105.000 110.800 105.500 112.100 ;
        RECT 107.800 110.800 108.200 113.100 ;
        RECT 109.400 110.800 109.800 112.100 ;
        RECT 111.600 110.800 112.000 113.500 ;
        RECT 114.200 110.800 114.600 113.300 ;
        RECT 116.600 110.800 117.000 113.000 ;
        RECT 119.400 110.800 119.800 112.100 ;
        RECT 121.000 110.800 121.500 112.100 ;
        RECT 123.800 110.800 124.200 113.100 ;
        RECT 125.400 110.800 125.800 113.100 ;
        RECT 127.000 110.800 127.400 113.100 ;
        RECT 128.600 110.800 129.000 113.100 ;
        RECT 130.200 110.800 130.600 113.100 ;
        RECT 131.800 110.800 132.200 113.100 ;
        RECT 133.400 110.800 133.800 113.300 ;
        RECT 136.000 110.800 136.400 113.500 ;
        RECT 138.200 110.800 138.600 112.100 ;
        RECT 141.400 110.800 141.800 113.000 ;
        RECT 144.200 110.800 144.600 112.100 ;
        RECT 145.800 110.800 146.300 112.100 ;
        RECT 148.600 110.800 149.000 113.100 ;
        RECT 151.000 110.800 151.400 112.100 ;
        RECT 152.600 110.800 153.000 113.100 ;
        RECT 155.300 110.800 155.800 112.100 ;
        RECT 157.000 110.800 157.400 112.100 ;
        RECT 159.800 110.800 160.200 113.000 ;
        RECT 162.200 110.800 162.600 113.300 ;
        RECT 164.800 110.800 165.200 113.500 ;
        RECT 167.000 110.800 167.400 112.100 ;
        RECT 167.800 110.800 168.200 113.100 ;
        RECT 171.000 110.800 171.400 112.700 ;
        RECT 174.200 110.800 174.600 112.100 ;
        RECT 175.800 110.800 176.200 111.900 ;
        RECT 0.200 110.200 180.600 110.800 ;
        RECT 1.400 107.900 1.800 110.200 ;
        RECT 4.100 108.900 4.600 110.200 ;
        RECT 5.800 108.900 6.200 110.200 ;
        RECT 8.600 108.000 9.000 110.200 ;
        RECT 10.500 107.900 10.900 110.200 ;
        RECT 12.600 108.900 13.000 110.200 ;
        RECT 13.400 108.900 13.800 110.200 ;
        RECT 15.000 108.900 15.400 110.200 ;
        RECT 16.600 107.900 17.000 110.200 ;
        RECT 19.300 108.900 19.800 110.200 ;
        RECT 21.000 108.900 21.400 110.200 ;
        RECT 23.800 108.000 24.200 110.200 ;
        RECT 25.600 107.900 26.000 110.200 ;
        RECT 28.600 107.900 29.000 110.200 ;
        RECT 30.200 107.900 30.600 110.200 ;
        RECT 32.900 108.900 33.400 110.200 ;
        RECT 34.600 108.900 35.000 110.200 ;
        RECT 37.400 108.000 37.800 110.200 ;
        RECT 41.400 107.700 41.800 110.200 ;
        RECT 44.000 107.500 44.400 110.200 ;
        RECT 46.200 108.900 46.600 110.200 ;
        RECT 47.000 107.900 47.400 110.200 ;
        RECT 51.800 106.900 52.200 110.200 ;
        RECT 52.600 107.900 53.000 110.200 ;
        RECT 55.600 107.900 56.000 110.200 ;
        RECT 56.600 108.900 57.000 110.200 ;
        RECT 58.200 108.900 58.600 110.200 ;
        RECT 59.000 108.900 59.400 110.200 ;
        RECT 61.100 107.900 61.500 110.200 ;
        RECT 62.200 106.900 62.600 110.200 ;
        RECT 67.000 107.900 67.400 110.200 ;
        RECT 68.600 108.000 69.000 110.200 ;
        RECT 71.400 108.900 71.800 110.200 ;
        RECT 73.000 108.900 73.500 110.200 ;
        RECT 75.800 107.900 76.200 110.200 ;
        RECT 78.200 108.900 78.600 110.200 ;
        RECT 79.800 109.100 80.200 110.200 ;
        RECT 84.000 107.900 84.400 110.200 ;
        RECT 87.000 107.900 87.400 110.200 ;
        RECT 89.400 107.900 89.800 110.200 ;
        RECT 91.800 107.900 92.200 110.200 ;
        RECT 93.400 107.900 93.800 110.200 ;
        RECT 95.000 107.900 95.400 110.200 ;
        RECT 96.600 107.900 97.000 110.200 ;
        RECT 98.200 107.900 98.600 110.200 ;
        RECT 99.200 107.900 99.600 110.200 ;
        RECT 102.200 107.900 102.600 110.200 ;
        RECT 103.000 107.900 103.400 110.200 ;
        RECT 104.600 107.900 105.000 110.200 ;
        RECT 105.600 107.900 106.000 110.200 ;
        RECT 108.600 107.900 109.000 110.200 ;
        RECT 109.400 108.900 109.800 110.200 ;
        RECT 111.800 108.000 112.200 110.200 ;
        RECT 114.600 108.900 115.000 110.200 ;
        RECT 116.200 108.900 116.700 110.200 ;
        RECT 119.000 107.900 119.400 110.200 ;
        RECT 121.400 107.900 121.800 110.200 ;
        RECT 124.100 108.900 124.600 110.200 ;
        RECT 125.800 108.900 126.200 110.200 ;
        RECT 128.600 108.000 129.000 110.200 ;
        RECT 131.000 107.900 131.400 110.200 ;
        RECT 133.700 108.900 134.200 110.200 ;
        RECT 135.400 108.900 135.800 110.200 ;
        RECT 138.200 108.000 138.600 110.200 ;
        RECT 141.400 108.900 141.800 110.200 ;
        RECT 143.600 107.500 144.000 110.200 ;
        RECT 146.200 107.700 146.600 110.200 ;
        RECT 147.800 108.900 148.200 110.200 ;
        RECT 150.200 108.000 150.600 110.200 ;
        RECT 153.000 108.900 153.400 110.200 ;
        RECT 154.600 108.900 155.100 110.200 ;
        RECT 157.400 107.900 157.800 110.200 ;
        RECT 159.800 108.300 160.200 110.200 ;
        RECT 163.000 108.300 163.400 110.200 ;
        RECT 166.500 107.900 166.900 110.200 ;
        RECT 168.600 108.900 169.000 110.200 ;
        RECT 170.200 108.900 170.600 110.200 ;
        RECT 171.800 108.000 172.200 110.200 ;
        RECT 174.600 108.900 175.000 110.200 ;
        RECT 176.200 108.900 176.700 110.200 ;
        RECT 179.000 107.900 179.400 110.200 ;
        RECT 1.400 90.800 1.800 93.100 ;
        RECT 4.100 90.800 4.600 92.100 ;
        RECT 5.800 90.800 6.200 92.100 ;
        RECT 8.600 90.800 9.000 93.000 ;
        RECT 10.200 90.800 10.600 92.100 ;
        RECT 12.400 90.800 12.800 93.500 ;
        RECT 15.000 90.800 15.400 93.300 ;
        RECT 16.800 90.800 17.200 93.100 ;
        RECT 19.800 90.800 20.200 93.100 ;
        RECT 20.600 90.800 21.000 92.100 ;
        RECT 22.200 90.800 22.600 92.100 ;
        RECT 23.000 90.800 23.400 92.100 ;
        RECT 25.100 90.800 25.500 93.100 ;
        RECT 27.000 90.800 27.400 93.000 ;
        RECT 29.800 90.800 30.200 92.100 ;
        RECT 31.400 90.800 31.900 92.100 ;
        RECT 34.200 90.800 34.600 93.100 ;
        RECT 35.800 90.800 36.200 94.100 ;
        RECT 41.900 90.800 42.300 93.000 ;
        RECT 46.200 90.800 46.600 94.100 ;
        RECT 47.000 90.800 47.400 94.100 ;
        RECT 51.800 90.800 52.200 93.100 ;
        RECT 55.800 90.800 56.200 91.900 ;
        RECT 57.400 90.800 57.800 92.100 ;
        RECT 59.800 90.800 60.200 93.100 ;
        RECT 62.500 90.800 63.000 92.100 ;
        RECT 64.200 90.800 64.600 92.100 ;
        RECT 67.000 90.800 67.400 93.000 ;
        RECT 68.600 90.800 69.000 92.100 ;
        RECT 70.800 90.800 71.200 93.500 ;
        RECT 73.400 90.800 73.800 93.300 ;
        RECT 75.800 90.800 76.200 93.000 ;
        RECT 78.600 90.800 79.000 92.100 ;
        RECT 80.200 90.800 80.700 92.100 ;
        RECT 83.000 90.800 83.400 93.100 ;
        RECT 87.000 90.800 87.400 93.000 ;
        RECT 89.800 90.800 90.200 92.100 ;
        RECT 91.400 90.800 91.900 92.100 ;
        RECT 94.200 90.800 94.600 93.100 ;
        RECT 95.800 90.800 96.200 93.100 ;
        RECT 98.200 90.800 98.600 93.100 ;
        RECT 101.400 90.800 101.800 93.000 ;
        RECT 104.200 90.800 104.600 92.100 ;
        RECT 105.800 90.800 106.300 92.100 ;
        RECT 108.600 90.800 109.000 93.100 ;
        RECT 110.800 90.800 111.200 93.500 ;
        RECT 113.400 90.800 113.800 93.300 ;
        RECT 115.000 90.800 115.400 92.100 ;
        RECT 116.600 90.800 117.000 92.100 ;
        RECT 117.400 90.800 117.800 92.100 ;
        RECT 120.600 90.800 121.000 93.100 ;
        RECT 126.200 90.800 126.600 92.100 ;
        RECT 127.800 90.800 128.200 92.100 ;
        RECT 132.600 90.800 133.000 93.100 ;
        RECT 138.200 90.800 138.600 93.100 ;
        RECT 143.000 90.800 143.400 92.100 ;
        RECT 144.600 90.800 145.000 92.100 ;
        RECT 150.200 90.800 150.600 93.100 ;
        RECT 153.400 90.800 153.800 92.100 ;
        RECT 154.800 90.800 155.200 93.500 ;
        RECT 157.400 90.800 157.800 93.300 ;
        RECT 159.600 90.800 160.000 93.500 ;
        RECT 162.200 90.800 162.600 93.300 ;
        RECT 164.600 90.800 165.000 92.100 ;
        RECT 166.200 90.800 166.600 93.000 ;
        RECT 169.000 90.800 169.400 92.100 ;
        RECT 170.600 90.800 171.100 92.100 ;
        RECT 173.400 90.800 173.800 93.100 ;
        RECT 175.800 90.800 176.200 93.100 ;
        RECT 178.200 90.800 178.600 93.100 ;
        RECT 0.200 90.200 180.600 90.800 ;
        RECT 1.400 87.900 1.800 90.200 ;
        RECT 4.100 88.900 4.600 90.200 ;
        RECT 5.800 88.900 6.200 90.200 ;
        RECT 8.600 88.000 9.000 90.200 ;
        RECT 10.200 88.900 10.600 90.200 ;
        RECT 12.300 87.900 12.700 90.200 ;
        RECT 13.400 88.900 13.800 90.200 ;
        RECT 15.000 88.900 15.400 90.200 ;
        RECT 15.800 87.900 16.200 90.200 ;
        RECT 19.300 88.000 19.700 90.200 ;
        RECT 21.400 87.900 21.800 90.200 ;
        RECT 26.200 86.900 26.600 90.200 ;
        RECT 28.600 87.900 29.000 90.200 ;
        RECT 30.200 88.900 30.600 90.200 ;
        RECT 31.800 89.100 32.200 90.200 ;
        RECT 35.800 86.900 36.200 90.200 ;
        RECT 40.600 87.900 41.000 90.200 ;
        RECT 43.600 87.900 44.000 90.200 ;
        RECT 44.600 87.900 45.000 90.200 ;
        RECT 47.800 88.000 48.200 90.200 ;
        RECT 50.600 88.900 51.000 90.200 ;
        RECT 52.200 88.900 52.700 90.200 ;
        RECT 55.000 87.900 55.400 90.200 ;
        RECT 56.900 87.900 57.300 90.200 ;
        RECT 59.000 88.900 59.400 90.200 ;
        RECT 59.800 88.900 60.200 90.200 ;
        RECT 61.400 88.900 61.800 90.200 ;
        RECT 62.200 87.900 62.600 90.200 ;
        RECT 67.000 86.900 67.400 90.200 ;
        RECT 67.800 87.900 68.200 90.200 ;
        RECT 70.200 88.900 70.600 90.200 ;
        RECT 71.800 88.900 72.200 90.200 ;
        RECT 72.600 88.900 73.000 90.200 ;
        RECT 74.700 87.900 75.100 90.200 ;
        RECT 76.600 87.700 77.000 90.200 ;
        RECT 79.200 87.500 79.600 90.200 ;
        RECT 82.200 87.900 82.600 90.200 ;
        RECT 83.000 87.900 83.400 90.200 ;
        RECT 85.400 88.900 85.800 90.200 ;
        RECT 89.200 87.500 89.600 90.200 ;
        RECT 91.800 87.700 92.200 90.200 ;
        RECT 93.400 88.900 93.800 90.200 ;
        RECT 95.000 88.900 95.400 90.200 ;
        RECT 95.800 88.900 96.200 90.200 ;
        RECT 97.900 87.900 98.300 90.200 ;
        RECT 99.600 87.500 100.000 90.200 ;
        RECT 102.200 87.700 102.600 90.200 ;
        RECT 104.600 87.900 105.000 90.200 ;
        RECT 107.300 88.900 107.800 90.200 ;
        RECT 109.000 88.900 109.400 90.200 ;
        RECT 111.800 88.000 112.200 90.200 ;
        RECT 113.400 88.900 113.800 90.200 ;
        RECT 115.000 88.900 115.400 90.200 ;
        RECT 117.100 87.900 117.500 90.200 ;
        RECT 118.800 87.500 119.200 90.200 ;
        RECT 121.400 87.700 121.800 90.200 ;
        RECT 123.800 88.900 124.200 90.200 ;
        RECT 125.400 87.900 125.800 90.200 ;
        RECT 128.100 88.900 128.600 90.200 ;
        RECT 129.800 88.900 130.200 90.200 ;
        RECT 132.600 88.000 133.000 90.200 ;
        RECT 134.500 87.900 134.900 90.200 ;
        RECT 136.600 88.900 137.000 90.200 ;
        RECT 137.400 88.900 137.800 90.200 ;
        RECT 139.000 88.900 139.400 90.200 ;
        RECT 143.000 87.900 143.400 90.200 ;
        RECT 147.800 88.900 148.200 90.200 ;
        RECT 149.400 88.900 149.800 90.200 ;
        RECT 155.000 87.900 155.400 90.200 ;
        RECT 158.200 88.900 158.600 90.200 ;
        RECT 159.300 87.900 159.700 90.200 ;
        RECT 161.400 88.900 161.800 90.200 ;
        RECT 162.200 88.900 162.600 90.200 ;
        RECT 163.800 88.900 164.200 90.200 ;
        RECT 165.400 88.300 165.800 90.200 ;
        RECT 169.400 88.300 169.800 90.200 ;
        RECT 172.600 88.900 173.000 90.200 ;
        RECT 174.200 89.100 174.600 90.200 ;
        RECT 179.000 87.900 179.400 90.200 ;
        RECT 1.400 70.800 1.800 73.100 ;
        RECT 4.100 70.800 4.600 72.100 ;
        RECT 5.800 70.800 6.200 72.100 ;
        RECT 8.600 70.800 9.000 73.000 ;
        RECT 11.000 70.800 11.400 72.100 ;
        RECT 11.800 70.800 12.200 73.100 ;
        RECT 14.200 70.800 14.600 72.100 ;
        RECT 16.400 70.800 16.800 73.500 ;
        RECT 19.000 70.800 19.400 73.300 ;
        RECT 20.600 70.800 21.000 73.100 ;
        RECT 23.000 70.800 23.400 74.100 ;
        RECT 27.000 70.800 27.400 73.100 ;
        RECT 29.700 70.800 30.200 72.100 ;
        RECT 31.400 70.800 31.800 72.100 ;
        RECT 34.200 70.800 34.600 73.000 ;
        RECT 35.800 70.800 36.200 72.100 ;
        RECT 39.600 70.800 40.000 73.500 ;
        RECT 42.200 70.800 42.600 73.300 ;
        RECT 43.800 70.800 44.200 73.100 ;
        RECT 47.000 70.800 47.400 73.100 ;
        RECT 49.700 70.800 50.200 72.100 ;
        RECT 51.400 70.800 51.800 72.100 ;
        RECT 54.200 70.800 54.600 73.000 ;
        RECT 57.400 70.800 57.800 73.100 ;
        RECT 59.000 70.800 59.400 73.000 ;
        RECT 61.800 70.800 62.200 72.100 ;
        RECT 63.400 70.800 63.900 72.100 ;
        RECT 66.200 70.800 66.600 73.100 ;
        RECT 67.800 70.800 68.200 72.100 ;
        RECT 70.000 70.800 70.400 73.500 ;
        RECT 72.600 70.800 73.000 73.300 ;
        RECT 76.600 70.800 77.000 74.100 ;
        RECT 78.200 70.800 78.600 73.100 ;
        RECT 79.800 70.800 80.200 72.100 ;
        RECT 80.800 70.800 81.200 73.100 ;
        RECT 83.800 70.800 84.200 73.100 ;
        RECT 87.000 70.800 87.400 73.000 ;
        RECT 89.800 70.800 90.200 72.100 ;
        RECT 91.400 70.800 91.900 72.100 ;
        RECT 94.200 70.800 94.600 73.100 ;
        RECT 95.800 70.800 96.200 73.100 ;
        RECT 98.200 70.800 98.600 73.100 ;
        RECT 99.800 70.800 100.200 73.100 ;
        RECT 100.600 70.800 101.000 72.100 ;
        RECT 102.200 70.800 102.600 72.100 ;
        RECT 103.000 70.800 103.400 72.100 ;
        RECT 104.600 70.800 105.000 72.100 ;
        RECT 106.200 70.800 106.600 73.300 ;
        RECT 108.800 70.800 109.200 73.500 ;
        RECT 111.000 70.800 111.400 72.700 ;
        RECT 114.200 70.800 114.600 72.100 ;
        RECT 118.200 70.800 118.600 71.900 ;
        RECT 119.800 70.800 120.200 72.100 ;
        RECT 123.800 70.800 124.200 72.700 ;
        RECT 126.200 70.800 126.600 73.300 ;
        RECT 128.800 70.800 129.200 73.500 ;
        RECT 131.000 70.800 131.400 72.100 ;
        RECT 132.400 70.800 132.800 73.500 ;
        RECT 135.000 70.800 135.400 73.300 ;
        RECT 139.000 70.800 139.400 73.000 ;
        RECT 141.800 70.800 142.200 72.100 ;
        RECT 143.400 70.800 143.900 72.100 ;
        RECT 146.200 70.800 146.600 73.100 ;
        RECT 149.400 70.800 149.800 73.100 ;
        RECT 154.200 70.800 154.600 72.100 ;
        RECT 155.800 70.800 156.200 72.100 ;
        RECT 161.400 70.800 161.800 73.100 ;
        RECT 164.600 70.800 165.000 72.100 ;
        RECT 166.200 70.800 166.600 73.300 ;
        RECT 168.800 70.800 169.200 73.500 ;
        RECT 171.000 70.800 171.400 73.000 ;
        RECT 173.800 70.800 174.200 72.100 ;
        RECT 175.400 70.800 175.900 72.100 ;
        RECT 178.200 70.800 178.600 73.100 ;
        RECT 0.200 70.200 180.600 70.800 ;
        RECT 0.600 67.900 1.000 70.200 ;
        RECT 2.200 67.900 2.600 70.200 ;
        RECT 3.800 67.900 4.200 70.200 ;
        RECT 5.400 67.700 5.800 70.200 ;
        RECT 8.000 67.500 8.400 70.200 ;
        RECT 10.200 68.000 10.600 70.200 ;
        RECT 13.000 68.900 13.400 70.200 ;
        RECT 14.600 68.900 15.100 70.200 ;
        RECT 17.400 67.900 17.800 70.200 ;
        RECT 19.800 67.700 20.200 70.200 ;
        RECT 22.400 67.500 22.800 70.200 ;
        RECT 25.400 67.900 25.800 70.200 ;
        RECT 27.000 68.900 27.400 70.200 ;
        RECT 28.600 68.000 29.000 70.200 ;
        RECT 31.400 68.900 31.800 70.200 ;
        RECT 33.000 68.900 33.500 70.200 ;
        RECT 35.800 67.900 36.200 70.200 ;
        RECT 39.800 68.000 40.200 70.200 ;
        RECT 42.600 68.900 43.000 70.200 ;
        RECT 44.200 68.900 44.700 70.200 ;
        RECT 47.000 67.900 47.400 70.200 ;
        RECT 48.900 67.900 49.300 70.200 ;
        RECT 51.000 68.900 51.400 70.200 ;
        RECT 51.800 68.900 52.200 70.200 ;
        RECT 53.400 68.900 53.800 70.200 ;
        RECT 55.000 68.900 55.400 70.200 ;
        RECT 56.600 69.100 57.000 70.200 ;
        RECT 60.600 68.900 61.000 70.200 ;
        RECT 62.200 68.900 62.600 70.200 ;
        RECT 63.000 68.900 63.400 70.200 ;
        RECT 65.100 67.900 65.500 70.200 ;
        RECT 66.200 67.900 66.600 70.200 ;
        RECT 67.800 67.900 68.200 70.200 ;
        RECT 68.600 67.900 69.000 70.200 ;
        RECT 71.000 67.900 71.400 70.200 ;
        RECT 73.700 68.900 74.200 70.200 ;
        RECT 75.400 68.900 75.800 70.200 ;
        RECT 78.200 68.000 78.600 70.200 ;
        RECT 79.800 68.900 80.200 70.200 ;
        RECT 82.000 67.500 82.400 70.200 ;
        RECT 84.600 67.700 85.000 70.200 ;
        RECT 86.200 67.900 86.600 70.200 ;
        RECT 89.200 67.900 89.600 70.200 ;
        RECT 92.600 68.000 93.000 70.200 ;
        RECT 95.400 68.900 95.800 70.200 ;
        RECT 97.000 68.900 97.500 70.200 ;
        RECT 99.800 67.900 100.200 70.200 ;
        RECT 101.400 68.900 101.800 70.200 ;
        RECT 103.600 67.500 104.000 70.200 ;
        RECT 106.200 67.700 106.600 70.200 ;
        RECT 108.600 67.900 109.000 70.200 ;
        RECT 111.300 68.900 111.800 70.200 ;
        RECT 113.000 68.900 113.400 70.200 ;
        RECT 115.800 68.000 116.200 70.200 ;
        RECT 117.400 68.900 117.800 70.200 ;
        RECT 119.000 68.900 119.400 70.200 ;
        RECT 120.600 67.700 121.000 70.200 ;
        RECT 123.200 67.500 123.600 70.200 ;
        RECT 125.400 67.900 125.800 70.200 ;
        RECT 128.100 68.900 128.600 70.200 ;
        RECT 129.800 68.900 130.200 70.200 ;
        RECT 132.600 68.000 133.000 70.200 ;
        RECT 134.200 68.900 134.600 70.200 ;
        RECT 138.200 68.300 138.600 70.200 ;
        RECT 143.800 68.300 144.200 70.200 ;
        RECT 146.200 68.900 146.600 70.200 ;
        RECT 147.800 69.100 148.200 70.200 ;
        RECT 152.100 67.900 152.500 70.200 ;
        RECT 154.200 68.900 154.600 70.200 ;
        RECT 156.600 68.300 157.000 70.200 ;
        RECT 158.800 67.500 159.200 70.200 ;
        RECT 161.400 67.700 161.800 70.200 ;
        RECT 165.400 68.300 165.800 70.200 ;
        RECT 167.000 68.900 167.400 70.200 ;
        RECT 168.600 68.900 169.000 70.200 ;
        RECT 170.200 68.000 170.600 70.200 ;
        RECT 173.000 68.900 173.400 70.200 ;
        RECT 174.600 68.900 175.100 70.200 ;
        RECT 177.400 67.900 177.800 70.200 ;
        RECT 179.000 68.900 179.400 70.200 ;
        RECT 1.200 50.800 1.600 53.500 ;
        RECT 3.800 50.800 4.200 53.300 ;
        RECT 6.200 50.800 6.600 52.100 ;
        RECT 7.000 50.800 7.400 53.100 ;
        RECT 10.000 50.800 10.400 53.100 ;
        RECT 11.800 50.800 12.200 53.100 ;
        RECT 14.500 50.800 15.000 52.100 ;
        RECT 16.200 50.800 16.600 52.100 ;
        RECT 19.000 50.800 19.400 53.000 ;
        RECT 22.200 50.800 22.600 53.100 ;
        RECT 23.000 50.800 23.400 53.100 ;
        RECT 25.700 50.800 26.100 53.100 ;
        RECT 27.800 50.800 28.200 52.100 ;
        RECT 28.600 50.800 29.000 52.100 ;
        RECT 30.200 50.800 30.600 52.100 ;
        RECT 31.800 50.800 32.200 53.100 ;
        RECT 34.500 50.800 35.000 52.100 ;
        RECT 36.200 50.800 36.600 52.100 ;
        RECT 39.000 50.800 39.400 53.000 ;
        RECT 42.400 50.800 42.800 53.100 ;
        RECT 45.400 50.800 45.800 53.100 ;
        RECT 48.600 50.800 49.000 54.100 ;
        RECT 51.000 50.800 51.400 53.100 ;
        RECT 51.800 50.800 52.200 53.100 ;
        RECT 53.400 50.800 53.800 53.100 ;
        RECT 54.200 50.800 54.600 52.100 ;
        RECT 55.800 50.800 56.200 52.100 ;
        RECT 57.400 50.800 57.800 53.000 ;
        RECT 60.200 50.800 60.600 52.100 ;
        RECT 61.800 50.800 62.300 52.100 ;
        RECT 64.600 50.800 65.000 53.100 ;
        RECT 66.200 50.800 66.600 52.100 ;
        RECT 67.800 50.800 68.200 52.100 ;
        RECT 68.600 50.800 69.000 52.100 ;
        RECT 70.200 50.800 70.600 52.100 ;
        RECT 71.000 50.800 71.400 52.100 ;
        RECT 72.600 50.800 73.000 52.100 ;
        RECT 74.200 50.800 74.600 53.300 ;
        RECT 76.800 50.800 77.200 53.500 ;
        RECT 79.000 50.800 79.400 52.100 ;
        RECT 80.000 50.800 80.400 53.100 ;
        RECT 83.000 50.800 83.400 53.100 ;
        RECT 84.600 50.800 85.000 53.000 ;
        RECT 87.400 50.800 87.800 52.100 ;
        RECT 89.000 50.800 89.500 52.100 ;
        RECT 91.800 50.800 92.200 53.100 ;
        RECT 95.300 50.800 95.700 53.100 ;
        RECT 97.400 50.800 97.800 52.100 ;
        RECT 98.200 50.800 98.600 52.100 ;
        RECT 99.800 50.800 100.200 52.100 ;
        RECT 101.400 50.800 101.800 53.000 ;
        RECT 104.200 50.800 104.600 52.100 ;
        RECT 105.800 50.800 106.300 52.100 ;
        RECT 108.600 50.800 109.000 53.100 ;
        RECT 110.200 50.800 110.600 52.100 ;
        RECT 112.400 50.800 112.800 53.500 ;
        RECT 115.000 50.800 115.400 53.300 ;
        RECT 116.600 50.800 117.000 52.100 ;
        RECT 118.200 50.800 118.600 53.100 ;
        RECT 119.800 50.800 120.200 53.100 ;
        RECT 123.800 50.800 124.200 51.900 ;
        RECT 125.400 50.800 125.800 52.100 ;
        RECT 127.800 50.800 128.200 53.000 ;
        RECT 130.600 50.800 131.000 52.100 ;
        RECT 132.200 50.800 132.700 52.100 ;
        RECT 135.000 50.800 135.400 53.100 ;
        RECT 136.600 50.800 137.000 52.100 ;
        RECT 140.400 50.800 140.800 53.500 ;
        RECT 143.000 50.800 143.400 53.300 ;
        RECT 145.400 50.800 145.800 53.100 ;
        RECT 148.100 50.800 148.600 52.100 ;
        RECT 149.800 50.800 150.200 52.100 ;
        RECT 152.600 50.800 153.000 53.000 ;
        RECT 155.000 50.800 155.400 53.300 ;
        RECT 157.600 50.800 158.000 53.500 ;
        RECT 159.800 50.800 160.200 52.100 ;
        RECT 161.400 50.800 161.800 51.900 ;
        RECT 166.200 50.800 166.600 53.300 ;
        RECT 168.800 50.800 169.200 53.500 ;
        RECT 171.000 50.800 171.400 53.000 ;
        RECT 173.800 50.800 174.200 52.100 ;
        RECT 175.400 50.800 175.900 52.100 ;
        RECT 178.200 50.800 178.600 53.100 ;
        RECT 0.200 50.200 180.600 50.800 ;
        RECT 1.400 47.900 1.800 50.200 ;
        RECT 4.100 48.900 4.600 50.200 ;
        RECT 5.800 48.900 6.200 50.200 ;
        RECT 8.600 48.000 9.000 50.200 ;
        RECT 10.200 48.900 10.600 50.200 ;
        RECT 12.400 47.500 12.800 50.200 ;
        RECT 15.000 47.700 15.400 50.200 ;
        RECT 17.400 48.900 17.800 50.200 ;
        RECT 18.200 47.900 18.600 50.200 ;
        RECT 20.600 47.900 21.000 50.200 ;
        RECT 22.200 47.900 22.600 50.200 ;
        RECT 23.800 47.900 24.200 50.200 ;
        RECT 25.400 47.900 25.800 50.200 ;
        RECT 27.000 47.900 27.400 50.200 ;
        RECT 28.600 47.700 29.000 50.200 ;
        RECT 31.200 47.500 31.600 50.200 ;
        RECT 33.400 48.900 33.800 50.200 ;
        RECT 36.600 47.900 37.000 50.200 ;
        RECT 39.300 48.900 39.800 50.200 ;
        RECT 41.000 48.900 41.400 50.200 ;
        RECT 43.800 48.000 44.200 50.200 ;
        RECT 45.400 47.900 45.800 50.200 ;
        RECT 47.000 47.900 47.400 50.200 ;
        RECT 48.600 47.900 49.000 50.200 ;
        RECT 50.200 47.900 50.600 50.200 ;
        RECT 51.800 47.900 52.200 50.200 ;
        RECT 52.600 48.900 53.000 50.200 ;
        RECT 54.200 48.900 54.600 50.200 ;
        RECT 55.000 48.900 55.400 50.200 ;
        RECT 57.100 47.900 57.500 50.200 ;
        RECT 58.200 48.900 58.600 50.200 ;
        RECT 59.800 48.900 60.200 50.200 ;
        RECT 63.800 49.100 64.200 50.200 ;
        RECT 65.400 48.900 65.800 50.200 ;
        RECT 67.000 47.900 67.400 50.200 ;
        RECT 70.200 48.900 70.600 50.200 ;
        RECT 71.800 47.900 72.200 50.200 ;
        RECT 74.500 48.900 75.000 50.200 ;
        RECT 76.200 48.900 76.600 50.200 ;
        RECT 79.000 48.000 79.400 50.200 ;
        RECT 81.400 47.900 81.800 50.200 ;
        RECT 84.100 48.900 84.600 50.200 ;
        RECT 85.800 48.900 86.200 50.200 ;
        RECT 88.600 48.000 89.000 50.200 ;
        RECT 92.600 47.700 93.000 50.200 ;
        RECT 95.200 47.500 95.600 50.200 ;
        RECT 97.400 48.900 97.800 50.200 ;
        RECT 98.400 47.900 98.800 50.200 ;
        RECT 101.400 47.900 101.800 50.200 ;
        RECT 102.400 47.900 102.800 50.200 ;
        RECT 105.400 47.900 105.800 50.200 ;
        RECT 106.200 47.900 106.600 50.200 ;
        RECT 107.800 48.900 108.200 50.200 ;
        RECT 110.200 47.900 110.600 50.200 ;
        RECT 112.900 48.900 113.400 50.200 ;
        RECT 114.600 48.900 115.000 50.200 ;
        RECT 117.400 48.000 117.800 50.200 ;
        RECT 120.600 48.300 121.000 50.200 ;
        RECT 122.200 48.900 122.600 50.200 ;
        RECT 124.600 48.300 125.000 50.200 ;
        RECT 127.600 47.500 128.000 50.200 ;
        RECT 130.200 47.700 130.600 50.200 ;
        RECT 131.800 48.900 132.200 50.200 ;
        RECT 134.200 47.700 134.600 50.200 ;
        RECT 136.800 47.500 137.200 50.200 ;
        RECT 139.000 48.900 139.400 50.200 ;
        RECT 141.400 47.900 141.800 50.200 ;
        RECT 143.000 47.900 143.400 50.200 ;
        RECT 144.600 47.900 145.000 50.200 ;
        RECT 146.200 47.900 146.600 50.200 ;
        RECT 147.800 47.900 148.200 50.200 ;
        RECT 149.400 47.700 149.800 50.200 ;
        RECT 152.000 47.500 152.400 50.200 ;
        RECT 154.200 48.300 154.600 50.200 ;
        RECT 157.400 48.000 157.800 50.200 ;
        RECT 160.200 48.900 160.600 50.200 ;
        RECT 161.800 48.900 162.300 50.200 ;
        RECT 164.600 47.900 165.000 50.200 ;
        RECT 167.000 48.300 167.400 50.200 ;
        RECT 170.200 48.900 170.600 50.200 ;
        RECT 171.800 48.000 172.200 50.200 ;
        RECT 174.600 48.900 175.000 50.200 ;
        RECT 176.200 48.900 176.700 50.200 ;
        RECT 179.000 47.900 179.400 50.200 ;
        RECT 1.400 30.800 1.800 33.100 ;
        RECT 4.100 30.800 4.600 32.100 ;
        RECT 5.800 30.800 6.200 32.100 ;
        RECT 8.600 30.800 9.000 33.000 ;
        RECT 10.800 30.800 11.200 33.500 ;
        RECT 13.400 30.800 13.800 33.300 ;
        RECT 15.200 30.800 15.600 33.100 ;
        RECT 18.200 30.800 18.600 33.100 ;
        RECT 19.800 30.800 20.200 33.100 ;
        RECT 22.500 30.800 23.000 32.100 ;
        RECT 24.200 30.800 24.600 32.100 ;
        RECT 27.000 30.800 27.400 33.000 ;
        RECT 29.400 30.800 29.800 33.300 ;
        RECT 32.000 30.800 32.400 33.500 ;
        RECT 34.200 30.800 34.600 32.100 ;
        RECT 35.800 30.800 36.200 33.300 ;
        RECT 38.400 30.800 38.800 33.500 ;
        RECT 42.200 30.800 42.600 32.100 ;
        RECT 45.400 30.800 45.800 34.100 ;
        RECT 46.200 30.800 46.600 34.100 ;
        RECT 49.400 30.800 49.800 34.100 ;
        RECT 53.400 30.800 53.800 33.100 ;
        RECT 54.200 30.800 54.600 34.100 ;
        RECT 57.400 30.800 57.800 32.100 ;
        RECT 59.000 30.800 59.400 32.100 ;
        RECT 60.600 30.800 61.000 32.900 ;
        RECT 62.200 30.800 62.600 32.100 ;
        RECT 63.000 30.800 63.400 32.100 ;
        RECT 64.600 30.800 65.000 33.100 ;
        RECT 67.800 30.800 68.200 32.100 ;
        RECT 69.400 30.800 69.800 31.900 ;
        RECT 75.000 30.800 75.400 33.100 ;
        RECT 75.800 30.800 76.200 32.100 ;
        RECT 77.400 30.800 77.800 32.100 ;
        RECT 78.200 30.800 78.600 32.100 ;
        RECT 79.800 30.800 80.200 32.100 ;
        RECT 80.600 30.800 81.000 32.100 ;
        RECT 82.200 30.800 82.600 32.100 ;
        RECT 83.000 30.800 83.400 33.100 ;
        RECT 86.000 30.800 86.400 33.100 ;
        RECT 89.400 30.800 89.800 33.300 ;
        RECT 92.000 30.800 92.400 33.500 ;
        RECT 94.200 30.800 94.600 32.100 ;
        RECT 95.800 30.800 96.200 33.100 ;
        RECT 98.500 30.800 99.000 32.100 ;
        RECT 100.200 30.800 100.600 32.100 ;
        RECT 103.000 30.800 103.400 33.000 ;
        RECT 104.600 30.800 105.000 32.100 ;
        RECT 106.200 30.800 106.600 32.100 ;
        RECT 107.000 30.800 107.400 32.100 ;
        RECT 109.100 30.800 109.500 33.100 ;
        RECT 111.000 30.800 111.400 33.000 ;
        RECT 113.800 30.800 114.200 32.100 ;
        RECT 115.400 30.800 115.900 32.100 ;
        RECT 118.200 30.800 118.600 33.100 ;
        RECT 120.600 30.800 121.000 32.700 ;
        RECT 123.000 30.800 123.400 32.100 ;
        RECT 124.600 30.800 125.000 32.900 ;
        RECT 126.200 30.800 126.600 33.100 ;
        RECT 127.800 30.800 128.200 33.100 ;
        RECT 129.400 30.800 129.800 33.100 ;
        RECT 131.000 30.800 131.400 33.100 ;
        RECT 132.600 30.800 133.000 33.100 ;
        RECT 134.200 30.800 134.600 33.100 ;
        RECT 136.900 30.800 137.400 32.100 ;
        RECT 138.600 30.800 139.000 32.100 ;
        RECT 141.400 30.800 141.800 33.000 ;
        RECT 146.200 30.800 146.600 32.700 ;
        RECT 148.600 30.800 149.000 33.100 ;
        RECT 151.300 30.800 151.800 32.100 ;
        RECT 153.000 30.800 153.400 32.100 ;
        RECT 155.800 30.800 156.200 33.000 ;
        RECT 157.400 30.800 157.800 32.100 ;
        RECT 159.000 30.800 159.400 32.100 ;
        RECT 161.200 30.800 161.600 33.500 ;
        RECT 163.800 30.800 164.200 33.300 ;
        RECT 166.200 30.800 166.600 33.000 ;
        RECT 169.000 30.800 169.400 32.100 ;
        RECT 170.600 30.800 171.100 32.100 ;
        RECT 173.400 30.800 173.800 33.100 ;
        RECT 175.800 30.800 176.200 33.300 ;
        RECT 178.400 30.800 178.800 33.500 ;
        RECT 0.200 30.200 180.600 30.800 ;
        RECT 1.400 27.900 1.800 30.200 ;
        RECT 4.100 28.900 4.600 30.200 ;
        RECT 5.800 28.900 6.200 30.200 ;
        RECT 8.600 28.000 9.000 30.200 ;
        RECT 10.200 28.900 10.600 30.200 ;
        RECT 12.400 27.500 12.800 30.200 ;
        RECT 15.000 27.700 15.400 30.200 ;
        RECT 16.800 27.900 17.200 30.200 ;
        RECT 19.800 27.900 20.200 30.200 ;
        RECT 20.600 27.900 21.000 30.200 ;
        RECT 22.200 27.900 22.600 30.200 ;
        RECT 23.800 27.900 24.200 30.200 ;
        RECT 25.400 27.900 25.800 30.200 ;
        RECT 27.000 27.900 27.400 30.200 ;
        RECT 28.600 27.900 29.000 30.200 ;
        RECT 31.300 28.900 31.800 30.200 ;
        RECT 33.000 28.900 33.400 30.200 ;
        RECT 35.800 28.000 36.200 30.200 ;
        RECT 39.000 27.900 39.400 30.200 ;
        RECT 41.400 27.900 41.800 30.200 ;
        RECT 44.400 27.900 44.800 30.200 ;
        RECT 47.000 27.900 47.400 30.200 ;
        RECT 50.200 26.900 50.600 30.200 ;
        RECT 51.000 26.900 51.400 30.200 ;
        RECT 55.000 27.900 55.400 30.200 ;
        RECT 55.800 27.900 56.200 30.200 ;
        RECT 59.000 28.900 59.400 30.200 ;
        RECT 59.800 27.900 60.200 30.200 ;
        RECT 62.200 28.900 62.600 30.200 ;
        RECT 63.800 28.900 64.200 30.200 ;
        RECT 66.200 27.900 66.600 30.200 ;
        RECT 67.800 28.900 68.200 30.200 ;
        RECT 69.400 28.100 69.800 30.200 ;
        RECT 71.000 28.900 71.400 30.200 ;
        RECT 75.000 29.100 75.400 30.200 ;
        RECT 76.600 28.900 77.000 30.200 ;
        RECT 78.200 27.900 78.600 30.200 ;
        RECT 81.400 28.900 81.800 30.200 ;
        RECT 83.000 28.000 83.400 30.200 ;
        RECT 85.800 28.900 86.200 30.200 ;
        RECT 87.400 28.900 87.900 30.200 ;
        RECT 90.200 27.900 90.600 30.200 ;
        RECT 93.400 28.900 93.800 30.200 ;
        RECT 95.600 27.500 96.000 30.200 ;
        RECT 98.200 27.700 98.600 30.200 ;
        RECT 100.600 27.700 101.000 30.200 ;
        RECT 103.200 27.500 103.600 30.200 ;
        RECT 105.400 28.900 105.800 30.200 ;
        RECT 107.000 28.000 107.400 30.200 ;
        RECT 109.800 28.900 110.200 30.200 ;
        RECT 111.400 28.900 111.900 30.200 ;
        RECT 114.200 27.900 114.600 30.200 ;
        RECT 117.400 27.900 117.800 30.200 ;
        RECT 119.000 27.700 119.400 30.200 ;
        RECT 121.600 27.500 122.000 30.200 ;
        RECT 123.800 28.900 124.200 30.200 ;
        RECT 126.200 27.900 126.600 30.200 ;
        RECT 127.800 28.000 128.200 30.200 ;
        RECT 130.600 28.900 131.000 30.200 ;
        RECT 132.200 28.900 132.700 30.200 ;
        RECT 135.000 27.900 135.400 30.200 ;
        RECT 138.200 28.300 138.600 30.200 ;
        RECT 143.000 27.900 143.400 30.200 ;
        RECT 143.800 28.900 144.200 30.200 ;
        RECT 146.200 28.000 146.600 30.200 ;
        RECT 149.000 28.900 149.400 30.200 ;
        RECT 150.600 28.900 151.100 30.200 ;
        RECT 153.400 27.900 153.800 30.200 ;
        RECT 155.000 28.900 155.400 30.200 ;
        RECT 158.200 27.900 158.600 30.200 ;
        RECT 159.800 28.900 160.200 30.200 ;
        RECT 161.400 27.900 161.800 30.200 ;
        RECT 164.100 28.900 164.600 30.200 ;
        RECT 165.800 28.900 166.200 30.200 ;
        RECT 168.600 28.000 169.000 30.200 ;
        RECT 171.000 28.900 171.400 30.200 ;
        RECT 173.400 28.300 173.800 30.200 ;
        RECT 175.800 28.300 176.200 30.200 ;
        RECT 179.800 27.900 180.200 30.200 ;
        RECT 1.200 10.800 1.600 13.500 ;
        RECT 3.800 10.800 4.200 13.300 ;
        RECT 6.200 10.800 6.600 12.100 ;
        RECT 7.300 10.800 7.700 13.100 ;
        RECT 9.400 10.800 9.800 12.100 ;
        RECT 10.200 10.800 10.600 12.100 ;
        RECT 11.800 10.800 12.200 12.100 ;
        RECT 13.400 10.800 13.800 13.000 ;
        RECT 16.200 10.800 16.600 12.100 ;
        RECT 17.800 10.800 18.300 12.100 ;
        RECT 20.600 10.800 21.000 13.100 ;
        RECT 23.000 10.800 23.400 13.300 ;
        RECT 25.600 10.800 26.000 13.500 ;
        RECT 27.800 10.800 28.200 12.100 ;
        RECT 29.400 10.800 29.800 13.100 ;
        RECT 32.100 10.800 32.600 12.100 ;
        RECT 33.800 10.800 34.200 12.100 ;
        RECT 36.600 10.800 37.000 13.000 ;
        RECT 40.600 10.800 41.000 13.300 ;
        RECT 43.200 10.800 43.600 13.500 ;
        RECT 44.600 10.800 45.000 12.100 ;
        RECT 47.000 10.800 47.400 13.000 ;
        RECT 49.800 10.800 50.200 12.100 ;
        RECT 51.400 10.800 51.900 12.100 ;
        RECT 54.200 10.800 54.600 13.100 ;
        RECT 55.800 10.800 56.200 12.100 ;
        RECT 57.400 10.800 57.800 12.100 ;
        RECT 58.200 10.800 58.600 12.100 ;
        RECT 60.300 10.800 60.700 13.100 ;
        RECT 61.400 10.800 61.800 12.100 ;
        RECT 63.600 10.800 64.000 13.500 ;
        RECT 66.200 10.800 66.600 13.300 ;
        RECT 69.400 10.800 69.800 13.100 ;
        RECT 70.200 10.800 70.600 12.100 ;
        RECT 71.800 10.800 72.200 12.100 ;
        RECT 72.600 10.800 73.000 12.100 ;
        RECT 74.700 10.800 75.100 13.100 ;
        RECT 75.800 10.800 76.200 13.100 ;
        RECT 77.400 10.800 77.800 13.100 ;
        RECT 79.000 10.800 79.400 13.100 ;
        RECT 80.600 10.800 81.000 13.000 ;
        RECT 83.400 10.800 83.800 12.100 ;
        RECT 85.000 10.800 85.500 12.100 ;
        RECT 87.800 10.800 88.200 13.100 ;
        RECT 91.000 10.800 91.400 12.100 ;
        RECT 93.200 10.800 93.600 13.500 ;
        RECT 95.800 10.800 96.200 13.300 ;
        RECT 98.200 10.800 98.600 13.000 ;
        RECT 101.000 10.800 101.400 12.100 ;
        RECT 102.600 10.800 103.100 12.100 ;
        RECT 105.400 10.800 105.800 13.100 ;
        RECT 107.000 10.800 107.400 12.100 ;
        RECT 109.200 10.800 109.600 13.500 ;
        RECT 111.800 10.800 112.200 13.300 ;
        RECT 113.400 10.800 113.800 12.100 ;
        RECT 115.800 10.800 116.200 13.300 ;
        RECT 118.400 10.800 118.800 13.500 ;
        RECT 119.800 10.800 120.200 12.100 ;
        RECT 122.200 10.800 122.600 13.300 ;
        RECT 124.800 10.800 125.200 13.500 ;
        RECT 127.000 10.800 127.400 13.100 ;
        RECT 129.700 10.800 130.200 12.100 ;
        RECT 131.400 10.800 131.800 12.100 ;
        RECT 134.200 10.800 134.600 13.000 ;
        RECT 135.800 10.800 136.200 12.100 ;
        RECT 138.000 10.800 138.400 13.500 ;
        RECT 140.600 10.800 141.000 13.300 ;
        RECT 144.400 10.800 144.800 13.500 ;
        RECT 147.000 10.800 147.400 13.300 ;
        RECT 149.400 10.800 149.800 13.300 ;
        RECT 152.000 10.800 152.400 13.500 ;
        RECT 154.200 10.800 154.600 13.100 ;
        RECT 156.900 10.800 157.400 12.100 ;
        RECT 158.600 10.800 159.000 12.100 ;
        RECT 161.400 10.800 161.800 13.000 ;
        RECT 163.800 10.800 164.200 13.300 ;
        RECT 166.400 10.800 166.800 13.500 ;
        RECT 167.800 10.800 168.200 13.100 ;
        RECT 171.000 10.800 171.400 12.100 ;
        RECT 171.800 10.800 172.200 12.100 ;
        RECT 174.200 10.800 174.600 12.100 ;
        RECT 175.600 10.800 176.000 13.500 ;
        RECT 178.200 10.800 178.600 13.300 ;
        RECT 0.200 10.200 180.600 10.800 ;
        RECT 1.400 7.900 1.800 10.200 ;
        RECT 4.100 8.900 4.600 10.200 ;
        RECT 5.800 8.900 6.200 10.200 ;
        RECT 8.600 8.000 9.000 10.200 ;
        RECT 11.000 7.900 11.400 10.200 ;
        RECT 13.700 8.900 14.200 10.200 ;
        RECT 15.400 8.900 15.800 10.200 ;
        RECT 18.200 8.000 18.600 10.200 ;
        RECT 20.100 7.900 20.500 10.200 ;
        RECT 22.200 8.900 22.600 10.200 ;
        RECT 23.000 8.900 23.400 10.200 ;
        RECT 24.600 8.900 25.000 10.200 ;
        RECT 26.200 7.900 26.600 10.200 ;
        RECT 28.900 8.900 29.400 10.200 ;
        RECT 30.600 8.900 31.000 10.200 ;
        RECT 33.400 8.000 33.800 10.200 ;
        RECT 37.400 7.900 37.800 10.200 ;
        RECT 40.100 8.900 40.600 10.200 ;
        RECT 41.800 8.900 42.200 10.200 ;
        RECT 44.600 8.000 45.000 10.200 ;
        RECT 46.200 8.900 46.600 10.200 ;
        RECT 47.800 8.900 48.200 10.200 ;
        RECT 48.600 8.900 49.000 10.200 ;
        RECT 50.700 7.900 51.100 10.200 ;
        RECT 52.600 7.900 53.000 10.200 ;
        RECT 55.300 8.900 55.800 10.200 ;
        RECT 57.000 8.900 57.400 10.200 ;
        RECT 59.800 8.000 60.200 10.200 ;
        RECT 61.400 7.900 61.800 10.200 ;
        RECT 63.000 7.900 63.400 10.200 ;
        RECT 64.600 7.900 65.000 10.200 ;
        RECT 66.200 8.000 66.600 10.200 ;
        RECT 69.000 8.900 69.400 10.200 ;
        RECT 70.600 8.900 71.100 10.200 ;
        RECT 73.400 7.900 73.800 10.200 ;
        RECT 75.800 7.900 76.200 10.200 ;
        RECT 78.500 8.900 79.000 10.200 ;
        RECT 80.200 8.900 80.600 10.200 ;
        RECT 83.000 8.000 83.400 10.200 ;
        RECT 84.600 8.900 85.000 10.200 ;
        RECT 86.800 7.500 87.200 10.200 ;
        RECT 89.400 7.700 89.800 10.200 ;
        RECT 92.600 7.900 93.000 10.200 ;
        RECT 94.200 7.900 94.600 10.200 ;
        RECT 95.800 7.900 96.200 10.200 ;
        RECT 97.400 8.000 97.800 10.200 ;
        RECT 100.200 8.900 100.600 10.200 ;
        RECT 101.800 8.900 102.300 10.200 ;
        RECT 104.600 7.900 105.000 10.200 ;
        RECT 107.800 7.900 108.200 10.200 ;
        RECT 109.400 7.900 109.800 10.200 ;
        RECT 112.100 8.900 112.600 10.200 ;
        RECT 113.800 8.900 114.200 10.200 ;
        RECT 116.600 8.000 117.000 10.200 ;
        RECT 118.200 7.900 118.600 10.200 ;
        RECT 119.800 7.900 120.200 10.200 ;
        RECT 121.400 7.900 121.800 10.200 ;
        RECT 122.200 8.900 122.600 10.200 ;
        RECT 123.800 8.900 124.200 10.200 ;
        RECT 125.400 8.900 125.800 10.200 ;
        RECT 127.000 7.900 127.400 10.200 ;
        RECT 129.700 8.900 130.200 10.200 ;
        RECT 131.400 8.900 131.800 10.200 ;
        RECT 134.200 8.000 134.600 10.200 ;
        RECT 135.800 7.900 136.200 10.200 ;
        RECT 138.200 8.900 138.600 10.200 ;
        RECT 142.000 7.500 142.400 10.200 ;
        RECT 144.600 7.700 145.000 10.200 ;
        RECT 147.000 7.700 147.400 10.200 ;
        RECT 149.600 7.500 150.000 10.200 ;
        RECT 151.800 7.900 152.200 10.200 ;
        RECT 154.500 8.900 155.000 10.200 ;
        RECT 156.200 8.900 156.600 10.200 ;
        RECT 159.000 8.000 159.400 10.200 ;
        RECT 161.400 7.900 161.800 10.200 ;
        RECT 164.100 8.900 164.600 10.200 ;
        RECT 165.800 8.900 166.200 10.200 ;
        RECT 168.600 8.000 169.000 10.200 ;
        RECT 171.000 7.900 171.400 10.200 ;
        RECT 173.700 8.900 174.200 10.200 ;
        RECT 175.400 8.900 175.800 10.200 ;
        RECT 178.200 8.000 178.600 10.200 ;
      LAYER via1 ;
        RECT 89.000 170.300 89.400 170.700 ;
        RECT 89.700 170.300 90.100 170.700 ;
        RECT 89.000 150.300 89.400 150.700 ;
        RECT 89.700 150.300 90.100 150.700 ;
        RECT 89.000 130.300 89.400 130.700 ;
        RECT 89.700 130.300 90.100 130.700 ;
        RECT 89.000 110.300 89.400 110.700 ;
        RECT 89.700 110.300 90.100 110.700 ;
        RECT 89.000 90.300 89.400 90.700 ;
        RECT 89.700 90.300 90.100 90.700 ;
        RECT 89.000 70.300 89.400 70.700 ;
        RECT 89.700 70.300 90.100 70.700 ;
        RECT 89.000 50.300 89.400 50.700 ;
        RECT 89.700 50.300 90.100 50.700 ;
        RECT 89.000 30.300 89.400 30.700 ;
        RECT 89.700 30.300 90.100 30.700 ;
        RECT 89.000 10.300 89.400 10.700 ;
        RECT 89.700 10.300 90.100 10.700 ;
      LAYER metal2 ;
        RECT 88.800 170.300 90.400 170.700 ;
        RECT 88.800 150.300 90.400 150.700 ;
        RECT 88.800 130.300 90.400 130.700 ;
        RECT 88.800 110.300 90.400 110.700 ;
        RECT 88.800 90.300 90.400 90.700 ;
        RECT 88.800 70.300 90.400 70.700 ;
        RECT 88.800 50.300 90.400 50.700 ;
        RECT 88.800 30.300 90.400 30.700 ;
        RECT 88.800 10.300 90.400 10.700 ;
      LAYER via2 ;
        RECT 89.000 170.300 89.400 170.700 ;
        RECT 89.700 170.300 90.100 170.700 ;
        RECT 89.000 150.300 89.400 150.700 ;
        RECT 89.700 150.300 90.100 150.700 ;
        RECT 89.000 130.300 89.400 130.700 ;
        RECT 89.700 130.300 90.100 130.700 ;
        RECT 89.000 110.300 89.400 110.700 ;
        RECT 89.700 110.300 90.100 110.700 ;
        RECT 89.000 90.300 89.400 90.700 ;
        RECT 89.700 90.300 90.100 90.700 ;
        RECT 89.000 70.300 89.400 70.700 ;
        RECT 89.700 70.300 90.100 70.700 ;
        RECT 89.000 50.300 89.400 50.700 ;
        RECT 89.700 50.300 90.100 50.700 ;
        RECT 89.000 30.300 89.400 30.700 ;
        RECT 89.700 30.300 90.100 30.700 ;
        RECT 89.000 10.300 89.400 10.700 ;
        RECT 89.700 10.300 90.100 10.700 ;
      LAYER metal3 ;
        RECT 88.800 170.300 90.400 170.700 ;
        RECT 88.800 150.300 90.400 150.700 ;
        RECT 88.800 130.300 90.400 130.700 ;
        RECT 88.800 110.300 90.400 110.700 ;
        RECT 88.800 90.300 90.400 90.700 ;
        RECT 88.800 70.300 90.400 70.700 ;
        RECT 88.800 50.300 90.400 50.700 ;
        RECT 88.800 30.300 90.400 30.700 ;
        RECT 88.800 10.300 90.400 10.700 ;
      LAYER via3 ;
        RECT 89.000 170.300 89.400 170.700 ;
        RECT 89.800 170.300 90.200 170.700 ;
        RECT 89.000 150.300 89.400 150.700 ;
        RECT 89.800 150.300 90.200 150.700 ;
        RECT 89.000 130.300 89.400 130.700 ;
        RECT 89.800 130.300 90.200 130.700 ;
        RECT 89.000 110.300 89.400 110.700 ;
        RECT 89.800 110.300 90.200 110.700 ;
        RECT 89.000 90.300 89.400 90.700 ;
        RECT 89.800 90.300 90.200 90.700 ;
        RECT 89.000 70.300 89.400 70.700 ;
        RECT 89.800 70.300 90.200 70.700 ;
        RECT 89.000 50.300 89.400 50.700 ;
        RECT 89.800 50.300 90.200 50.700 ;
        RECT 89.000 30.300 89.400 30.700 ;
        RECT 89.800 30.300 90.200 30.700 ;
        RECT 89.000 10.300 89.400 10.700 ;
        RECT 89.800 10.300 90.200 10.700 ;
      LAYER metal4 ;
        RECT 88.800 170.300 90.400 170.700 ;
        RECT 88.800 150.300 90.400 150.700 ;
        RECT 88.800 130.300 90.400 130.700 ;
        RECT 88.800 110.300 90.400 110.700 ;
        RECT 88.800 90.300 90.400 90.700 ;
        RECT 88.800 70.300 90.400 70.700 ;
        RECT 88.800 50.300 90.400 50.700 ;
        RECT 88.800 30.300 90.400 30.700 ;
        RECT 88.800 10.300 90.400 10.700 ;
      LAYER via4 ;
        RECT 89.000 170.300 89.400 170.700 ;
        RECT 89.700 170.300 90.100 170.700 ;
        RECT 89.000 150.300 89.400 150.700 ;
        RECT 89.700 150.300 90.100 150.700 ;
        RECT 89.000 130.300 89.400 130.700 ;
        RECT 89.700 130.300 90.100 130.700 ;
        RECT 89.000 110.300 89.400 110.700 ;
        RECT 89.700 110.300 90.100 110.700 ;
        RECT 89.000 90.300 89.400 90.700 ;
        RECT 89.700 90.300 90.100 90.700 ;
        RECT 89.000 70.300 89.400 70.700 ;
        RECT 89.700 70.300 90.100 70.700 ;
        RECT 89.000 50.300 89.400 50.700 ;
        RECT 89.700 50.300 90.100 50.700 ;
        RECT 89.000 30.300 89.400 30.700 ;
        RECT 89.700 30.300 90.100 30.700 ;
        RECT 89.000 10.300 89.400 10.700 ;
        RECT 89.700 10.300 90.100 10.700 ;
      LAYER metal5 ;
        RECT 88.800 170.200 90.400 170.700 ;
        RECT 88.800 150.200 90.400 150.700 ;
        RECT 88.800 130.200 90.400 130.700 ;
        RECT 88.800 110.200 90.400 110.700 ;
        RECT 88.800 90.200 90.400 90.700 ;
        RECT 88.800 70.200 90.400 70.700 ;
        RECT 88.800 50.200 90.400 50.700 ;
        RECT 88.800 30.200 90.400 30.700 ;
        RECT 88.800 10.200 90.400 10.700 ;
      LAYER via5 ;
        RECT 89.800 170.200 90.300 170.700 ;
        RECT 89.800 150.200 90.300 150.700 ;
        RECT 89.800 130.200 90.300 130.700 ;
        RECT 89.800 110.200 90.300 110.700 ;
        RECT 89.800 90.200 90.300 90.700 ;
        RECT 89.800 70.200 90.300 70.700 ;
        RECT 89.800 50.200 90.300 50.700 ;
        RECT 89.800 30.200 90.300 30.700 ;
        RECT 89.800 10.200 90.300 10.700 ;
      LAYER metal6 ;
        RECT 88.800 -3.000 90.400 173.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 59.800 166.900 60.200 167.200 ;
        RECT 59.300 166.500 60.200 166.900 ;
        RECT 74.200 166.900 74.600 167.200 ;
        RECT 74.200 166.500 75.100 166.900 ;
        RECT 33.700 154.100 34.600 154.500 ;
        RECT 34.200 153.800 34.600 154.100 ;
        RECT 147.000 154.100 147.900 154.500 ;
        RECT 147.000 153.800 147.400 154.100 ;
        RECT 131.300 114.100 132.200 114.500 ;
        RECT 131.800 113.800 132.200 114.100 ;
        RECT 98.200 106.900 98.600 107.200 ;
        RECT 97.700 106.500 98.600 106.900 ;
        RECT 27.000 46.900 27.400 47.200 ;
        RECT 26.500 46.500 27.400 46.900 ;
        RECT 45.400 46.900 45.800 47.200 ;
        RECT 147.800 46.900 148.200 47.200 ;
        RECT 45.400 46.500 46.300 46.900 ;
        RECT 147.300 46.500 148.200 46.900 ;
        RECT 132.100 34.100 133.000 34.500 ;
        RECT 132.600 33.800 133.000 34.100 ;
        RECT 27.000 26.900 27.400 27.200 ;
        RECT 26.500 26.500 27.400 26.900 ;
      LAYER via1 ;
        RECT 59.800 166.800 60.200 167.200 ;
        RECT 74.200 166.800 74.600 167.200 ;
        RECT 98.200 106.800 98.600 107.200 ;
        RECT 27.000 46.800 27.400 47.200 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 27.000 26.800 27.400 27.200 ;
      LAYER metal2 ;
        RECT 59.800 172.800 60.200 173.200 ;
        RECT 59.800 167.200 60.100 172.800 ;
        RECT 59.800 166.800 60.200 167.200 ;
        RECT 74.200 166.800 74.600 167.200 ;
        RECT 59.800 163.200 60.100 166.800 ;
        RECT 74.200 163.200 74.500 166.800 ;
        RECT 34.200 162.800 34.600 163.200 ;
        RECT 59.800 162.800 60.200 163.200 ;
        RECT 74.200 162.800 74.600 163.200 ;
        RECT 34.200 154.200 34.500 162.800 ;
        RECT 34.200 153.800 34.600 154.200 ;
        RECT 146.200 154.100 146.600 154.200 ;
        RECT 147.000 154.100 147.400 154.200 ;
        RECT 146.200 153.800 147.400 154.100 ;
        RECT 131.800 114.100 132.200 114.200 ;
        RECT 132.600 114.100 133.000 114.200 ;
        RECT 131.800 113.800 133.000 114.100 ;
        RECT 98.200 107.800 98.600 108.200 ;
        RECT 98.200 107.200 98.500 107.800 ;
        RECT 98.200 106.800 98.600 107.200 ;
        RECT 27.000 47.800 27.400 48.200 ;
        RECT 45.400 47.800 45.800 48.200 ;
        RECT 27.000 47.200 27.300 47.800 ;
        RECT 45.400 47.200 45.700 47.800 ;
        RECT 27.000 46.800 27.400 47.200 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 147.800 46.800 148.200 47.200 ;
        RECT 27.000 27.200 27.300 46.800 ;
        RECT 45.400 41.200 45.700 46.800 ;
        RECT 147.800 45.200 148.100 46.800 ;
        RECT 132.600 44.800 133.000 45.200 ;
        RECT 147.800 44.800 148.200 45.200 ;
        RECT 132.600 41.200 132.900 44.800 ;
        RECT 45.400 40.800 45.800 41.200 ;
        RECT 132.600 40.800 133.000 41.200 ;
        RECT 132.600 34.200 132.900 40.800 ;
        RECT 132.600 33.800 133.000 34.200 ;
        RECT 27.000 26.800 27.400 27.200 ;
      LAYER via2 ;
        RECT 132.600 113.800 133.000 114.200 ;
      LAYER metal3 ;
        RECT 34.200 163.100 34.600 163.200 ;
        RECT 59.800 163.100 60.200 163.200 ;
        RECT 74.200 163.100 74.600 163.200 ;
        RECT 131.800 163.100 132.200 163.200 ;
        RECT 34.200 162.800 132.200 163.100 ;
        RECT 131.800 154.100 132.200 154.200 ;
        RECT 146.200 154.100 146.600 154.200 ;
        RECT 131.800 153.800 146.600 154.100 ;
        RECT 131.800 114.100 132.200 114.200 ;
        RECT 132.600 114.100 133.000 114.200 ;
        RECT 131.800 113.800 133.000 114.100 ;
        RECT 98.200 108.100 98.600 108.200 ;
        RECT 131.800 108.100 132.200 108.200 ;
        RECT 98.200 107.800 132.200 108.100 ;
        RECT 27.000 48.100 27.400 48.200 ;
        RECT 45.400 48.100 45.800 48.200 ;
        RECT 27.000 47.800 45.800 48.100 ;
        RECT 131.800 45.100 132.200 45.200 ;
        RECT 132.600 45.100 133.000 45.200 ;
        RECT 147.800 45.100 148.200 45.200 ;
        RECT 131.800 44.800 148.200 45.100 ;
        RECT 45.400 41.100 45.800 41.200 ;
        RECT 132.600 41.100 133.000 41.200 ;
        RECT 45.400 40.800 133.000 41.100 ;
      LAYER via3 ;
        RECT 131.800 162.800 132.200 163.200 ;
        RECT 131.800 107.800 132.200 108.200 ;
      LAYER metal4 ;
        RECT 131.800 162.800 132.200 163.200 ;
        RECT 131.800 154.200 132.100 162.800 ;
        RECT 131.800 153.800 132.200 154.200 ;
        RECT 131.800 114.200 132.100 153.800 ;
        RECT 131.800 113.800 132.200 114.200 ;
        RECT 131.800 108.200 132.100 113.800 ;
        RECT 131.800 107.800 132.200 108.200 ;
        RECT 131.800 45.200 132.100 107.800 ;
        RECT 131.800 44.800 132.200 45.200 ;
    END
  END clk
  PIN rst_n
    PORT
      LAYER metal1 ;
        RECT 121.400 166.000 121.800 166.300 ;
        RECT 130.200 166.000 130.600 166.200 ;
        RECT 131.800 166.000 132.200 166.200 ;
        RECT 136.600 166.100 136.900 166.200 ;
        RECT 132.700 166.000 133.100 166.100 ;
        RECT 121.400 165.700 133.100 166.000 ;
        RECT 136.500 166.000 136.900 166.100 ;
        RECT 139.000 166.000 139.400 166.200 ;
        RECT 147.800 166.000 148.200 166.300 ;
        RECT 136.500 165.700 148.200 166.000 ;
        RECT 136.600 165.200 136.900 165.700 ;
        RECT 136.600 164.800 137.000 165.200 ;
        RECT 156.500 155.000 168.200 155.300 ;
        RECT 156.500 154.900 156.900 155.000 ;
        RECT 157.400 154.800 157.800 155.000 ;
        RECT 159.000 154.800 159.400 155.000 ;
        RECT 167.800 154.700 168.200 155.000 ;
        RECT 162.900 146.000 163.300 146.100 ;
        RECT 164.600 146.000 165.000 146.200 ;
        RECT 165.400 146.000 165.800 146.200 ;
        RECT 174.200 146.000 174.600 146.300 ;
        RECT 162.900 145.700 174.600 146.000 ;
        RECT 122.200 95.000 133.900 95.300 ;
        RECT 122.200 94.700 122.600 95.000 ;
        RECT 131.000 94.800 131.400 95.000 ;
        RECT 132.600 94.800 133.000 95.000 ;
        RECT 133.500 94.900 133.900 95.000 ;
        RECT 137.300 95.000 149.000 95.300 ;
        RECT 137.300 94.900 137.800 95.000 ;
        RECT 137.400 94.800 137.800 94.900 ;
        RECT 139.800 94.800 140.200 95.000 ;
        RECT 148.600 94.700 149.000 95.000 ;
        RECT 142.100 86.000 142.500 86.100 ;
        RECT 144.600 86.000 145.000 86.200 ;
        RECT 153.400 86.000 153.800 86.300 ;
        RECT 142.100 85.700 153.800 86.000 ;
        RECT 148.500 75.000 160.200 75.300 ;
        RECT 148.500 74.900 148.900 75.000 ;
        RECT 151.000 74.800 151.400 75.000 ;
        RECT 154.200 74.800 154.600 75.000 ;
        RECT 159.800 74.700 160.200 75.000 ;
      LAYER via1 ;
        RECT 130.200 165.800 130.600 166.200 ;
        RECT 131.800 165.800 132.200 166.200 ;
        RECT 147.800 165.800 148.200 166.200 ;
        RECT 164.600 145.800 165.000 146.200 ;
        RECT 148.600 94.800 149.000 95.200 ;
        RECT 153.400 85.800 153.800 86.200 ;
      LAYER metal2 ;
        RECT 130.200 172.800 130.600 173.200 ;
        RECT 130.200 166.200 130.500 172.800 ;
        RECT 130.200 165.800 130.600 166.200 ;
        RECT 131.800 166.100 132.200 166.200 ;
        RECT 132.600 166.100 133.000 166.200 ;
        RECT 131.800 165.800 133.000 166.100 ;
        RECT 136.600 165.800 137.000 166.200 ;
        RECT 147.800 165.800 148.200 166.200 ;
        RECT 136.600 165.200 136.900 165.800 ;
        RECT 136.600 164.800 137.000 165.200 ;
        RECT 147.800 155.200 148.100 165.800 ;
        RECT 157.400 155.800 157.800 156.200 ;
        RECT 157.400 155.200 157.700 155.800 ;
        RECT 147.800 154.800 148.200 155.200 ;
        RECT 157.400 154.800 157.800 155.200 ;
        RECT 157.400 149.200 157.700 154.800 ;
        RECT 157.400 148.800 157.800 149.200 ;
        RECT 164.600 148.800 165.000 149.200 ;
        RECT 164.600 146.200 164.900 148.800 ;
        RECT 164.600 145.800 165.000 146.200 ;
        RECT 132.600 95.800 133.000 96.200 ;
        RECT 137.400 95.800 137.800 96.200 ;
        RECT 148.600 95.800 149.000 96.200 ;
        RECT 153.400 95.800 153.800 96.200 ;
        RECT 132.600 95.200 132.900 95.800 ;
        RECT 137.400 95.200 137.700 95.800 ;
        RECT 148.600 95.200 148.900 95.800 ;
        RECT 132.600 94.800 133.000 95.200 ;
        RECT 137.400 94.800 137.800 95.200 ;
        RECT 148.600 94.800 149.000 95.200 ;
        RECT 153.400 86.200 153.700 95.800 ;
        RECT 153.400 85.800 153.800 86.200 ;
        RECT 153.400 79.100 153.700 85.800 ;
        RECT 153.400 78.800 154.500 79.100 ;
        RECT 154.200 75.200 154.500 78.800 ;
        RECT 154.200 74.800 154.600 75.200 ;
      LAYER via2 ;
        RECT 132.600 165.800 133.000 166.200 ;
      LAYER metal3 ;
        RECT 132.600 166.100 133.000 166.200 ;
        RECT 136.600 166.100 137.000 166.200 ;
        RECT 132.600 165.800 137.000 166.100 ;
        RECT 157.400 155.800 157.800 156.200 ;
        RECT 147.800 155.100 148.200 155.200 ;
        RECT 148.600 155.100 149.000 155.200 ;
        RECT 157.400 155.100 157.700 155.800 ;
        RECT 147.800 154.800 157.700 155.100 ;
        RECT 157.400 149.100 157.800 149.200 ;
        RECT 164.600 149.100 165.000 149.200 ;
        RECT 157.400 148.800 165.000 149.100 ;
        RECT 148.600 96.800 149.000 97.200 ;
        RECT 148.600 96.200 148.900 96.800 ;
        RECT 132.600 96.100 133.000 96.200 ;
        RECT 137.400 96.100 137.800 96.200 ;
        RECT 132.600 95.800 137.800 96.100 ;
        RECT 148.600 96.100 149.000 96.200 ;
        RECT 153.400 96.100 153.800 96.200 ;
        RECT 148.600 95.800 153.800 96.100 ;
      LAYER via3 ;
        RECT 148.600 154.800 149.000 155.200 ;
      LAYER metal4 ;
        RECT 148.600 154.800 149.000 155.200 ;
        RECT 148.600 97.200 148.900 154.800 ;
        RECT 148.600 96.800 149.000 97.200 ;
    END
  END rst_n
  PIN cs
    PORT
      LAYER metal1 ;
        RECT 106.200 3.800 106.600 5.200 ;
      LAYER metal2 ;
        RECT 106.200 3.800 106.600 4.200 ;
        RECT 106.200 -1.900 106.500 3.800 ;
        RECT 107.000 -1.900 107.400 -1.800 ;
        RECT 106.200 -2.200 107.400 -1.900 ;
    END
  END cs
  PIN re
    PORT
      LAYER metal1 ;
        RECT 125.400 7.800 125.800 8.600 ;
      LAYER metal2 ;
        RECT 125.400 7.800 125.800 8.200 ;
        RECT 124.600 -1.900 125.000 -1.800 ;
        RECT 125.400 -1.900 125.700 7.800 ;
        RECT 124.600 -2.200 125.700 -1.900 ;
    END
  END re
  PIN we
    PORT
      LAYER metal1 ;
        RECT 122.200 7.800 122.600 8.600 ;
        RECT 107.800 6.800 108.200 7.600 ;
      LAYER metal2 ;
        RECT 122.200 8.100 122.600 8.200 ;
        RECT 123.000 8.100 123.400 8.200 ;
        RECT 122.200 7.800 123.400 8.100 ;
        RECT 107.800 6.800 108.200 7.200 ;
        RECT 107.800 4.200 108.100 6.800 ;
        RECT 107.800 3.800 108.200 4.200 ;
        RECT 107.800 -1.900 108.100 3.800 ;
        RECT 108.600 -1.900 109.000 -1.800 ;
        RECT 107.800 -2.200 109.000 -1.900 ;
      LAYER via2 ;
        RECT 123.000 7.800 123.400 8.200 ;
      LAYER metal3 ;
        RECT 122.200 8.100 122.600 8.200 ;
        RECT 123.000 8.100 123.400 8.200 ;
        RECT 122.200 7.800 123.400 8.100 ;
        RECT 107.800 4.100 108.200 4.200 ;
        RECT 122.200 4.100 122.600 4.200 ;
        RECT 107.800 3.800 122.600 4.100 ;
      LAYER via3 ;
        RECT 122.200 3.800 122.600 4.200 ;
      LAYER metal4 ;
        RECT 122.200 7.800 122.600 8.200 ;
        RECT 122.200 4.200 122.500 7.800 ;
        RECT 122.200 3.800 122.600 4.200 ;
    END
  END we
  PIN addr[0]
    PORT
      LAYER metal1 ;
        RECT 64.900 48.100 65.800 48.200 ;
        RECT 64.900 47.800 66.500 48.100 ;
        RECT 66.200 47.100 66.500 47.800 ;
        RECT 67.000 47.100 67.400 47.600 ;
        RECT 66.200 46.800 67.400 47.100 ;
        RECT 75.000 33.400 75.400 34.200 ;
        RECT 71.000 27.800 71.400 28.600 ;
        RECT 81.400 27.800 81.800 28.600 ;
      LAYER via1 ;
        RECT 67.000 46.800 67.400 47.200 ;
        RECT 75.000 33.800 75.400 34.200 ;
      LAYER metal2 ;
        RECT 67.000 46.800 67.400 47.200 ;
        RECT 67.000 37.200 67.300 46.800 ;
        RECT 67.000 36.800 67.400 37.200 ;
        RECT 71.000 36.800 71.400 37.200 ;
        RECT 75.000 36.800 75.400 37.200 ;
        RECT 71.000 28.200 71.300 36.800 ;
        RECT 75.000 34.200 75.300 36.800 ;
        RECT 75.000 33.800 75.400 34.200 ;
        RECT 71.000 27.800 71.400 28.200 ;
        RECT 80.600 28.100 81.000 28.200 ;
        RECT 81.400 28.100 81.800 28.200 ;
        RECT 80.600 27.800 81.800 28.100 ;
        RECT 81.400 14.100 81.700 27.800 ;
        RECT 80.600 13.800 81.700 14.100 ;
        RECT 80.600 -1.800 80.900 13.800 ;
        RECT 80.600 -2.200 81.000 -1.800 ;
      LAYER metal3 ;
        RECT 67.000 37.100 67.400 37.200 ;
        RECT 71.000 37.100 71.400 37.200 ;
        RECT 75.000 37.100 75.400 37.200 ;
        RECT 67.000 36.800 75.400 37.100 ;
        RECT 71.000 28.100 71.400 28.200 ;
        RECT 80.600 28.100 81.000 28.200 ;
        RECT 71.000 27.800 81.000 28.100 ;
    END
  END addr[0]
  PIN addr[1]
    PORT
      LAYER metal1 ;
        RECT 70.200 47.800 70.600 48.600 ;
        RECT 73.400 35.800 73.800 36.600 ;
        RECT 70.100 26.800 70.600 27.200 ;
        RECT 75.400 27.100 76.200 27.200 ;
        RECT 78.200 27.100 78.600 27.600 ;
        RECT 75.400 26.800 78.600 27.100 ;
        RECT 70.000 26.400 70.400 26.800 ;
      LAYER via1 ;
        RECT 70.200 26.800 70.600 27.200 ;
        RECT 75.800 26.800 76.200 27.200 ;
      LAYER metal2 ;
        RECT 70.200 47.800 70.600 48.200 ;
        RECT 70.200 36.200 70.500 47.800 ;
        RECT 70.200 35.800 70.600 36.200 ;
        RECT 72.600 36.100 73.000 36.200 ;
        RECT 73.400 36.100 73.800 36.200 ;
        RECT 72.600 35.800 73.800 36.100 ;
        RECT 70.200 27.200 70.500 35.800 ;
        RECT 70.200 26.800 70.600 27.200 ;
        RECT 75.000 27.100 75.400 27.200 ;
        RECT 75.800 27.100 76.200 27.200 ;
        RECT 75.000 26.800 76.200 27.100 ;
        RECT 70.200 -1.800 70.500 26.800 ;
        RECT 70.200 -2.200 70.600 -1.800 ;
      LAYER metal3 ;
        RECT 70.200 36.100 70.600 36.200 ;
        RECT 72.600 36.100 73.000 36.200 ;
        RECT 70.200 35.800 73.000 36.100 ;
        RECT 70.200 27.100 70.600 27.200 ;
        RECT 75.000 27.100 75.400 27.200 ;
        RECT 70.200 26.800 75.400 27.100 ;
    END
  END addr[1]
  PIN addr[2]
    PORT
      LAYER metal1 ;
        RECT 61.200 34.200 61.600 34.600 ;
        RECT 61.300 34.100 61.800 34.200 ;
        RECT 62.200 34.100 62.600 34.200 ;
        RECT 61.300 33.800 62.600 34.100 ;
        RECT 64.600 33.400 65.000 34.200 ;
        RECT 68.600 33.800 69.400 34.200 ;
        RECT 59.000 27.800 59.400 28.600 ;
        RECT 61.400 24.400 61.800 25.200 ;
      LAYER via1 ;
        RECT 62.200 33.800 62.600 34.200 ;
        RECT 64.600 33.800 65.000 34.200 ;
        RECT 61.400 24.800 61.800 25.200 ;
      LAYER metal2 ;
        RECT 68.600 34.800 69.000 35.200 ;
        RECT 68.600 34.200 68.900 34.800 ;
        RECT 62.200 34.100 62.600 34.200 ;
        RECT 63.000 34.100 63.400 34.200 ;
        RECT 62.200 33.800 63.400 34.100 ;
        RECT 63.800 34.100 64.200 34.200 ;
        RECT 64.600 34.100 65.000 34.200 ;
        RECT 63.800 33.800 65.000 34.100 ;
        RECT 68.600 33.800 69.000 34.200 ;
        RECT 63.000 30.200 63.300 33.800 ;
        RECT 59.000 29.800 59.400 30.200 ;
        RECT 63.000 29.800 63.400 30.200 ;
        RECT 59.000 28.200 59.300 29.800 ;
        RECT 59.000 27.800 59.400 28.200 ;
        RECT 63.000 26.200 63.300 29.800 ;
        RECT 61.400 25.800 61.800 26.200 ;
        RECT 62.200 25.800 62.600 26.200 ;
        RECT 63.000 25.800 63.400 26.200 ;
        RECT 61.400 25.200 61.700 25.800 ;
        RECT 61.400 24.800 61.800 25.200 ;
        RECT 61.400 -1.900 61.800 -1.800 ;
        RECT 62.200 -1.900 62.500 25.800 ;
        RECT 61.400 -2.200 62.500 -1.900 ;
      LAYER via2 ;
        RECT 63.000 33.800 63.400 34.200 ;
      LAYER metal3 ;
        RECT 68.600 34.800 69.000 35.200 ;
        RECT 63.000 34.100 63.400 34.200 ;
        RECT 63.800 34.100 64.200 34.200 ;
        RECT 68.600 34.100 68.900 34.800 ;
        RECT 63.000 33.800 68.900 34.100 ;
        RECT 59.000 30.100 59.400 30.200 ;
        RECT 63.000 30.100 63.400 30.200 ;
        RECT 59.000 29.800 63.400 30.100 ;
        RECT 61.400 26.100 61.800 26.200 ;
        RECT 62.200 26.100 62.600 26.200 ;
        RECT 63.000 26.100 63.400 26.200 ;
        RECT 61.400 25.800 63.400 26.100 ;
    END
  END addr[2]
  PIN addr[3]
    PORT
      LAYER metal1 ;
        RECT 62.200 33.100 62.600 33.200 ;
        RECT 63.000 33.100 63.400 33.200 ;
        RECT 62.200 32.800 63.400 33.100 ;
        RECT 62.200 32.400 62.600 32.800 ;
        RECT 63.000 32.400 63.400 32.800 ;
        RECT 55.800 26.800 56.200 27.600 ;
        RECT 59.800 26.800 60.200 27.600 ;
      LAYER metal2 ;
        RECT 62.200 32.800 62.600 33.200 ;
        RECT 62.200 28.200 62.500 32.800 ;
        RECT 59.800 27.800 60.200 28.200 ;
        RECT 62.200 27.800 62.600 28.200 ;
        RECT 59.800 27.200 60.100 27.800 ;
        RECT 55.800 26.800 56.200 27.200 ;
        RECT 59.800 26.800 60.200 27.200 ;
        RECT 55.800 26.200 56.100 26.800 ;
        RECT 59.800 26.200 60.100 26.800 ;
        RECT 55.800 25.800 56.200 26.200 ;
        RECT 59.800 25.800 60.200 26.200 ;
        RECT 56.600 0.800 57.000 1.200 ;
        RECT 56.600 -1.800 56.900 0.800 ;
        RECT 56.600 -2.200 57.000 -1.800 ;
      LAYER metal3 ;
        RECT 59.800 28.100 60.200 28.200 ;
        RECT 62.200 28.100 62.600 28.200 ;
        RECT 59.800 27.800 62.600 28.100 ;
        RECT 55.800 26.100 56.200 26.200 ;
        RECT 57.400 26.100 57.800 26.200 ;
        RECT 59.800 26.100 60.200 26.200 ;
        RECT 55.800 25.800 60.200 26.100 ;
        RECT 56.600 1.100 57.000 1.200 ;
        RECT 57.400 1.100 57.800 1.200 ;
        RECT 56.600 0.800 57.800 1.100 ;
      LAYER via3 ;
        RECT 57.400 25.800 57.800 26.200 ;
        RECT 57.400 0.800 57.800 1.200 ;
      LAYER metal4 ;
        RECT 57.400 25.800 57.800 26.200 ;
        RECT 57.400 1.200 57.700 25.800 ;
        RECT 57.400 0.800 57.800 1.200 ;
    END
  END addr[3]
  PIN din[0]
    PORT
      LAYER metal1 ;
        RECT 85.400 166.800 85.800 167.600 ;
      LAYER metal2 ;
        RECT 87.000 172.800 87.400 173.200 ;
        RECT 87.000 168.200 87.300 172.800 ;
        RECT 85.400 167.800 85.800 168.200 ;
        RECT 87.000 167.800 87.400 168.200 ;
        RECT 85.400 167.200 85.700 167.800 ;
        RECT 85.400 166.800 85.800 167.200 ;
      LAYER metal3 ;
        RECT 85.400 168.100 85.800 168.200 ;
        RECT 87.000 168.100 87.400 168.200 ;
        RECT 85.400 167.800 87.400 168.100 ;
    END
  END din[0]
  PIN din[1]
    PORT
      LAYER metal1 ;
        RECT 81.400 166.800 81.800 167.600 ;
      LAYER metal2 ;
        RECT 83.000 172.800 83.400 173.200 ;
        RECT 83.000 168.200 83.300 172.800 ;
        RECT 81.400 167.800 81.800 168.200 ;
        RECT 83.000 167.800 83.400 168.200 ;
        RECT 81.400 167.200 81.700 167.800 ;
        RECT 81.400 166.800 81.800 167.200 ;
      LAYER metal3 ;
        RECT 81.400 168.100 81.800 168.200 ;
        RECT 83.000 168.100 83.400 168.200 ;
        RECT 81.400 167.800 83.400 168.100 ;
    END
  END din[1]
  PIN din[2]
    PORT
      LAYER metal1 ;
        RECT 64.600 6.800 65.000 7.600 ;
      LAYER metal2 ;
        RECT 64.600 6.800 65.000 7.200 ;
        RECT 64.600 1.200 64.900 6.800 ;
        RECT 63.000 0.800 63.400 1.200 ;
        RECT 64.600 0.800 65.000 1.200 ;
        RECT 63.000 -1.800 63.300 0.800 ;
        RECT 63.000 -2.200 63.400 -1.800 ;
      LAYER metal3 ;
        RECT 63.000 1.100 63.400 1.200 ;
        RECT 64.600 1.100 65.000 1.200 ;
        RECT 63.000 0.800 65.000 1.100 ;
    END
  END din[2]
  PIN din[3]
    PORT
      LAYER metal1 ;
        RECT 70.200 166.800 70.600 167.600 ;
      LAYER metal2 ;
        RECT 71.800 172.800 72.200 173.200 ;
        RECT 71.800 168.200 72.100 172.800 ;
        RECT 70.200 167.800 70.600 168.200 ;
        RECT 71.800 167.800 72.200 168.200 ;
        RECT 70.200 167.200 70.500 167.800 ;
        RECT 70.200 166.800 70.600 167.200 ;
      LAYER metal3 ;
        RECT 70.200 168.100 70.600 168.200 ;
        RECT 71.800 168.100 72.200 168.200 ;
        RECT 70.200 167.800 72.200 168.100 ;
    END
  END din[3]
  PIN din[4]
    PORT
      LAYER metal1 ;
        RECT 79.000 13.400 79.400 14.200 ;
      LAYER via1 ;
        RECT 79.000 13.800 79.400 14.200 ;
      LAYER metal2 ;
        RECT 79.000 13.800 79.400 14.200 ;
        RECT 79.000 1.200 79.300 13.800 ;
        RECT 77.400 0.800 77.800 1.200 ;
        RECT 79.000 0.800 79.400 1.200 ;
        RECT 77.400 -1.800 77.700 0.800 ;
        RECT 77.400 -2.200 77.800 -1.800 ;
      LAYER metal3 ;
        RECT 77.400 1.100 77.800 1.200 ;
        RECT 79.000 1.100 79.400 1.200 ;
        RECT 77.400 0.800 79.400 1.100 ;
    END
  END din[4]
  PIN din[5]
    PORT
      LAYER metal1 ;
        RECT 121.400 6.800 121.800 7.600 ;
      LAYER metal2 ;
        RECT 119.800 7.800 120.200 8.200 ;
        RECT 121.400 7.800 121.800 8.200 ;
        RECT 119.800 -1.800 120.100 7.800 ;
        RECT 121.400 7.200 121.700 7.800 ;
        RECT 121.400 6.800 121.800 7.200 ;
        RECT 119.800 -2.200 120.200 -1.800 ;
      LAYER metal3 ;
        RECT 119.800 8.100 120.200 8.200 ;
        RECT 121.400 8.100 121.800 8.200 ;
        RECT 119.800 7.800 121.800 8.100 ;
    END
  END din[5]
  PIN din[6]
    PORT
      LAYER metal1 ;
        RECT 0.600 66.800 1.000 67.600 ;
      LAYER metal2 ;
        RECT 0.600 66.800 1.000 67.200 ;
        RECT 0.600 65.200 0.900 66.800 ;
        RECT 0.600 64.800 1.000 65.200 ;
      LAYER metal3 ;
        RECT -2.600 65.100 -2.200 65.200 ;
        RECT 0.600 65.100 1.000 65.200 ;
        RECT -2.600 64.800 1.000 65.100 ;
    END
  END din[6]
  PIN din[7]
    PORT
      LAYER metal1 ;
        RECT 95.800 6.800 96.200 7.600 ;
      LAYER metal2 ;
        RECT 95.800 6.800 96.200 7.200 ;
        RECT 95.800 1.200 96.100 6.800 ;
        RECT 94.200 0.800 94.600 1.200 ;
        RECT 95.800 0.800 96.200 1.200 ;
        RECT 94.200 -1.800 94.500 0.800 ;
        RECT 94.200 -2.200 94.600 -1.800 ;
      LAYER metal3 ;
        RECT 94.200 1.100 94.600 1.200 ;
        RECT 95.800 1.100 96.200 1.200 ;
        RECT 94.200 0.800 96.200 1.100 ;
    END
  END din[7]
  PIN dout[0]
    PORT
      LAYER metal1 ;
        RECT 155.000 166.200 155.400 169.900 ;
        RECT 155.100 165.100 155.400 166.200 ;
        RECT 155.000 161.100 155.400 165.100 ;
      LAYER via1 ;
        RECT 155.000 168.800 155.400 169.200 ;
      LAYER metal2 ;
        RECT 155.000 169.800 155.400 170.200 ;
        RECT 155.000 169.200 155.300 169.800 ;
        RECT 155.000 168.800 155.400 169.200 ;
      LAYER metal3 ;
        RECT 183.000 171.800 183.400 172.200 ;
        RECT 183.000 171.100 183.300 171.800 ;
        RECT 182.200 170.800 183.300 171.100 ;
        RECT 155.000 170.100 155.400 170.200 ;
        RECT 182.200 170.100 182.500 170.800 ;
        RECT 155.000 169.800 182.500 170.100 ;
    END
  END dout[0]
  PIN dout[1]
    PORT
      LAYER metal1 ;
        RECT 176.600 166.200 177.000 169.900 ;
        RECT 176.700 165.100 177.000 166.200 ;
        RECT 176.600 161.100 177.000 165.100 ;
      LAYER via1 ;
        RECT 176.600 168.800 177.000 169.200 ;
      LAYER metal2 ;
        RECT 176.600 168.800 177.000 169.200 ;
        RECT 176.600 168.200 176.900 168.800 ;
        RECT 176.600 167.800 177.000 168.200 ;
      LAYER metal3 ;
        RECT 183.000 169.800 183.400 170.200 ;
        RECT 183.000 169.100 183.300 169.800 ;
        RECT 176.600 168.800 183.300 169.100 ;
        RECT 176.600 168.200 176.900 168.800 ;
        RECT 176.600 167.800 177.000 168.200 ;
    END
  END dout[1]
  PIN dout[2]
    PORT
      LAYER metal1 ;
        RECT 175.000 155.900 175.400 159.900 ;
        RECT 175.100 154.800 175.400 155.900 ;
        RECT 175.000 151.100 175.400 154.800 ;
      LAYER via1 ;
        RECT 175.000 158.800 175.400 159.200 ;
      LAYER metal2 ;
        RECT 175.000 166.800 175.400 167.200 ;
        RECT 175.000 159.200 175.300 166.800 ;
        RECT 175.000 158.800 175.400 159.200 ;
      LAYER metal3 ;
        RECT 183.000 167.800 183.400 168.200 ;
        RECT 175.000 167.100 175.400 167.200 ;
        RECT 183.000 167.100 183.300 167.800 ;
        RECT 175.000 166.800 183.300 167.100 ;
    END
  END dout[2]
  PIN dout[3]
    PORT
      LAYER metal1 ;
        RECT 179.000 159.100 179.400 159.900 ;
        RECT 179.800 159.100 180.200 159.200 ;
        RECT 179.000 158.800 180.200 159.100 ;
        RECT 179.000 155.900 179.400 158.800 ;
        RECT 179.100 154.800 179.400 155.900 ;
        RECT 179.000 151.100 179.400 154.800 ;
      LAYER via1 ;
        RECT 179.800 158.800 180.200 159.200 ;
      LAYER metal2 ;
        RECT 179.800 165.800 180.200 166.200 ;
        RECT 179.800 159.200 180.100 165.800 ;
        RECT 179.800 158.800 180.200 159.200 ;
      LAYER metal3 ;
        RECT 179.800 166.100 180.200 166.200 ;
        RECT 183.000 166.100 183.400 166.200 ;
        RECT 179.800 165.800 183.400 166.100 ;
    END
  END dout[3]
  PIN dout[4]
    PORT
      LAYER metal1 ;
        RECT 176.600 95.900 177.000 99.900 ;
        RECT 176.700 94.800 177.000 95.900 ;
        RECT 176.600 91.100 177.000 94.800 ;
      LAYER via1 ;
        RECT 176.600 98.800 177.000 99.200 ;
      LAYER metal2 ;
        RECT 176.600 104.800 177.000 105.200 ;
        RECT 176.600 99.200 176.900 104.800 ;
        RECT 176.600 98.800 177.000 99.200 ;
      LAYER metal3 ;
        RECT 178.200 164.100 178.600 164.200 ;
        RECT 183.000 164.100 183.400 164.200 ;
        RECT 178.200 163.800 183.400 164.100 ;
        RECT 176.600 105.100 177.000 105.200 ;
        RECT 178.200 105.100 178.600 105.200 ;
        RECT 176.600 104.800 178.600 105.100 ;
      LAYER via3 ;
        RECT 178.200 104.800 178.600 105.200 ;
      LAYER metal4 ;
        RECT 178.200 163.800 178.600 164.200 ;
        RECT 178.200 105.200 178.500 163.800 ;
        RECT 178.200 104.800 178.600 105.200 ;
    END
  END dout[4]
  PIN dout[5]
    PORT
      LAYER metal1 ;
        RECT 179.000 95.900 179.400 99.900 ;
        RECT 179.100 94.800 179.400 95.900 ;
        RECT 179.000 91.100 179.400 94.800 ;
      LAYER via1 ;
        RECT 179.000 98.800 179.400 99.200 ;
      LAYER metal2 ;
        RECT 179.000 156.800 179.400 157.200 ;
        RECT 179.000 99.200 179.300 156.800 ;
        RECT 179.000 98.800 179.400 99.200 ;
      LAYER metal3 ;
        RECT 179.800 162.100 180.200 162.200 ;
        RECT 183.000 162.100 183.400 162.200 ;
        RECT 179.800 161.800 183.400 162.100 ;
        RECT 179.000 157.100 179.400 157.200 ;
        RECT 179.800 157.100 180.200 157.200 ;
        RECT 179.000 156.800 180.200 157.100 ;
      LAYER via3 ;
        RECT 179.800 156.800 180.200 157.200 ;
      LAYER metal4 ;
        RECT 179.800 161.800 180.200 162.200 ;
        RECT 179.800 157.200 180.100 161.800 ;
        RECT 179.800 156.800 180.200 157.200 ;
    END
  END dout[5]
  PIN dout[6]
    PORT
      LAYER metal1 ;
        RECT 179.800 86.200 180.200 89.900 ;
        RECT 179.900 85.100 180.200 86.200 ;
        RECT 179.800 81.100 180.200 85.100 ;
      LAYER via1 ;
        RECT 179.800 88.800 180.200 89.200 ;
      LAYER metal2 ;
        RECT 179.800 103.800 180.200 104.200 ;
        RECT 179.800 89.200 180.100 103.800 ;
        RECT 179.800 88.800 180.200 89.200 ;
      LAYER metal3 ;
        RECT 179.000 160.100 179.400 160.200 ;
        RECT 183.000 160.100 183.400 160.200 ;
        RECT 179.000 159.800 183.400 160.100 ;
        RECT 179.000 104.100 179.400 104.200 ;
        RECT 179.800 104.100 180.200 104.200 ;
        RECT 179.000 103.800 180.200 104.100 ;
      LAYER metal4 ;
        RECT 179.000 159.800 179.400 160.200 ;
        RECT 179.000 104.200 179.300 159.800 ;
        RECT 179.000 103.800 179.400 104.200 ;
    END
  END dout[6]
  PIN dout[7]
    PORT
      LAYER metal1 ;
        RECT 179.000 166.200 179.400 169.900 ;
        RECT 179.100 165.100 179.400 166.200 ;
        RECT 179.000 161.100 179.400 165.100 ;
      LAYER via1 ;
        RECT 179.000 161.800 179.400 162.200 ;
      LAYER metal2 ;
        RECT 179.000 161.800 179.400 162.200 ;
        RECT 179.000 158.200 179.300 161.800 ;
        RECT 179.000 157.800 179.400 158.200 ;
      LAYER metal3 ;
        RECT 179.000 158.100 179.400 158.200 ;
        RECT 183.000 158.100 183.400 158.200 ;
        RECT 179.000 157.800 183.400 158.100 ;
    END
  END dout[7]
  OBS
      LAYER metal1 ;
        RECT 0.600 166.100 1.000 169.900 ;
        RECT 1.400 167.800 1.800 168.600 ;
        RECT 4.100 168.000 4.500 169.500 ;
        RECT 6.200 168.500 6.600 169.500 ;
        RECT 3.700 167.700 4.500 168.000 ;
        RECT 3.700 167.500 4.100 167.700 ;
        RECT 3.700 167.200 4.000 167.500 ;
        RECT 6.300 167.400 6.600 168.500 ;
        RECT 7.000 167.500 7.400 169.900 ;
        RECT 9.200 169.200 9.600 169.900 ;
        RECT 8.600 168.900 9.600 169.200 ;
        RECT 11.400 168.900 11.800 169.900 ;
        RECT 13.500 169.200 14.100 169.900 ;
        RECT 13.400 168.900 14.100 169.200 ;
        RECT 8.600 168.500 9.000 168.900 ;
        RECT 11.400 168.600 11.700 168.900 ;
        RECT 9.400 168.200 9.800 168.600 ;
        RECT 10.300 168.300 11.700 168.600 ;
        RECT 13.400 168.500 13.800 168.900 ;
        RECT 10.300 168.200 10.700 168.300 ;
        RECT 3.000 166.800 4.000 167.200 ;
        RECT 4.500 167.100 6.600 167.400 ;
        RECT 7.400 167.100 8.200 167.200 ;
        RECT 9.500 167.100 9.800 168.200 ;
        RECT 14.300 167.700 14.700 167.800 ;
        RECT 15.800 167.700 16.200 169.900 ;
        RECT 14.300 167.400 16.200 167.700 ;
        RECT 16.600 167.500 17.000 169.900 ;
        RECT 18.800 169.200 19.200 169.900 ;
        RECT 18.200 168.900 19.200 169.200 ;
        RECT 21.000 168.900 21.400 169.900 ;
        RECT 23.100 169.200 23.700 169.900 ;
        RECT 23.000 168.900 23.700 169.200 ;
        RECT 18.200 168.500 18.600 168.900 ;
        RECT 21.000 168.600 21.300 168.900 ;
        RECT 19.000 168.200 19.400 168.600 ;
        RECT 19.900 168.300 21.300 168.600 ;
        RECT 23.000 168.500 23.400 168.900 ;
        RECT 19.900 168.200 20.300 168.300 ;
        RECT 12.300 167.100 12.700 167.200 ;
        RECT 4.500 166.900 5.000 167.100 ;
        RECT 3.000 166.100 3.400 166.200 ;
        RECT 0.600 165.800 3.400 166.100 ;
        RECT 0.600 161.100 1.000 165.800 ;
        RECT 3.000 165.400 3.400 165.800 ;
        RECT 3.700 165.200 4.000 166.800 ;
        RECT 4.300 166.500 5.000 166.900 ;
        RECT 7.400 166.800 12.900 167.100 ;
        RECT 8.900 166.700 9.300 166.800 ;
        RECT 4.700 165.500 5.000 166.500 ;
        RECT 5.400 165.800 5.800 166.600 ;
        RECT 6.200 165.800 6.600 166.600 ;
        RECT 8.100 166.200 8.500 166.300 ;
        RECT 9.400 166.200 9.800 166.300 ;
        RECT 12.600 166.200 12.900 166.800 ;
        RECT 13.400 166.400 13.800 166.500 ;
        RECT 8.100 165.900 10.600 166.200 ;
        RECT 10.200 165.800 10.600 165.900 ;
        RECT 12.600 165.800 13.000 166.200 ;
        RECT 13.400 166.100 15.300 166.400 ;
        RECT 14.900 166.000 15.300 166.100 ;
        RECT 7.000 165.500 9.800 165.600 ;
        RECT 4.700 165.200 6.600 165.500 ;
        RECT 3.700 164.900 4.200 165.200 ;
        RECT 3.700 164.600 4.500 164.900 ;
        RECT 4.100 161.100 4.500 164.600 ;
        RECT 6.300 163.500 6.600 165.200 ;
        RECT 6.200 161.500 6.600 163.500 ;
        RECT 7.000 165.400 9.900 165.500 ;
        RECT 7.000 165.300 11.900 165.400 ;
        RECT 7.000 161.100 7.400 165.300 ;
        RECT 9.500 165.100 11.900 165.300 ;
        RECT 8.600 164.500 11.300 164.800 ;
        RECT 8.600 164.400 9.000 164.500 ;
        RECT 10.900 164.400 11.300 164.500 ;
        RECT 11.600 164.500 11.900 165.100 ;
        RECT 12.600 165.200 12.900 165.800 ;
        RECT 14.100 165.700 14.500 165.800 ;
        RECT 15.800 165.700 16.200 167.400 ;
        RECT 17.000 167.100 17.800 167.200 ;
        RECT 19.100 167.100 19.400 168.200 ;
        RECT 23.900 167.700 24.300 167.800 ;
        RECT 25.400 167.700 25.800 169.900 ;
        RECT 23.900 167.400 25.800 167.700 ;
        RECT 21.900 167.100 22.300 167.200 ;
        RECT 17.000 166.800 22.500 167.100 ;
        RECT 18.500 166.700 18.900 166.800 ;
        RECT 17.700 166.200 18.100 166.300 ;
        RECT 22.200 166.200 22.500 166.800 ;
        RECT 23.000 166.400 23.400 166.500 ;
        RECT 17.700 166.100 20.200 166.200 ;
        RECT 20.600 166.100 21.000 166.200 ;
        RECT 17.700 165.900 21.000 166.100 ;
        RECT 19.800 165.800 21.000 165.900 ;
        RECT 22.200 165.800 22.600 166.200 ;
        RECT 23.000 166.100 24.900 166.400 ;
        RECT 24.500 166.000 24.900 166.100 ;
        RECT 14.100 165.400 16.200 165.700 ;
        RECT 12.600 164.900 13.800 165.200 ;
        RECT 12.300 164.500 12.700 164.600 ;
        RECT 11.600 164.200 12.700 164.500 ;
        RECT 13.500 164.400 13.800 164.900 ;
        RECT 13.500 164.000 14.200 164.400 ;
        RECT 10.300 163.700 10.700 163.800 ;
        RECT 11.700 163.700 12.100 163.800 ;
        RECT 8.600 163.100 9.000 163.500 ;
        RECT 10.300 163.400 12.100 163.700 ;
        RECT 11.400 163.100 11.700 163.400 ;
        RECT 13.400 163.100 13.800 163.500 ;
        RECT 8.600 162.800 9.600 163.100 ;
        RECT 9.200 161.100 9.600 162.800 ;
        RECT 11.400 161.100 11.800 163.100 ;
        RECT 13.500 161.100 14.100 163.100 ;
        RECT 15.800 161.100 16.200 165.400 ;
        RECT 16.600 165.500 19.400 165.600 ;
        RECT 16.600 165.400 19.500 165.500 ;
        RECT 16.600 165.300 21.500 165.400 ;
        RECT 16.600 161.100 17.000 165.300 ;
        RECT 19.100 165.100 21.500 165.300 ;
        RECT 18.200 164.500 20.900 164.800 ;
        RECT 18.200 164.400 18.600 164.500 ;
        RECT 20.500 164.400 20.900 164.500 ;
        RECT 21.200 164.500 21.500 165.100 ;
        RECT 22.200 165.200 22.500 165.800 ;
        RECT 23.700 165.700 24.100 165.800 ;
        RECT 25.400 165.700 25.800 167.400 ;
        RECT 23.700 165.400 25.800 165.700 ;
        RECT 22.200 164.900 23.400 165.200 ;
        RECT 21.900 164.500 22.300 164.600 ;
        RECT 21.200 164.200 22.300 164.500 ;
        RECT 23.100 164.400 23.400 164.900 ;
        RECT 23.100 164.000 23.800 164.400 ;
        RECT 19.900 163.700 20.300 163.800 ;
        RECT 21.300 163.700 21.700 163.800 ;
        RECT 18.200 163.100 18.600 163.500 ;
        RECT 19.900 163.400 21.700 163.700 ;
        RECT 21.000 163.100 21.300 163.400 ;
        RECT 23.000 163.100 23.400 163.500 ;
        RECT 18.200 162.800 19.200 163.100 ;
        RECT 18.800 161.100 19.200 162.800 ;
        RECT 21.000 161.100 21.400 163.100 ;
        RECT 23.100 161.100 23.700 163.100 ;
        RECT 25.400 161.100 25.800 165.400 ;
        RECT 26.200 167.700 26.600 169.900 ;
        RECT 28.300 169.200 28.900 169.900 ;
        RECT 28.300 168.900 29.000 169.200 ;
        RECT 30.600 168.900 31.000 169.900 ;
        RECT 32.800 169.200 33.200 169.900 ;
        RECT 32.800 168.900 33.800 169.200 ;
        RECT 28.600 168.500 29.000 168.900 ;
        RECT 30.700 168.600 31.000 168.900 ;
        RECT 30.700 168.300 32.100 168.600 ;
        RECT 31.700 168.200 32.100 168.300 ;
        RECT 32.600 168.200 33.000 168.600 ;
        RECT 33.400 168.500 33.800 168.900 ;
        RECT 27.700 167.700 28.100 167.800 ;
        RECT 26.200 167.400 28.100 167.700 ;
        RECT 26.200 165.700 26.600 167.400 ;
        RECT 29.700 167.100 30.100 167.200 ;
        RECT 32.600 167.100 32.900 168.200 ;
        RECT 35.000 167.500 35.400 169.900 ;
        RECT 37.400 168.500 37.800 169.500 ;
        RECT 37.400 167.400 37.700 168.500 ;
        RECT 39.500 168.000 39.900 169.500 ;
        RECT 39.500 167.700 40.300 168.000 ;
        RECT 39.900 167.500 40.300 167.700 ;
        RECT 34.200 167.100 35.000 167.200 ;
        RECT 37.400 167.100 39.500 167.400 ;
        RECT 29.500 166.800 35.000 167.100 ;
        RECT 39.000 166.900 39.500 167.100 ;
        RECT 40.000 167.200 40.300 167.500 ;
        RECT 40.000 167.100 41.000 167.200 ;
        RECT 41.400 167.100 41.800 167.200 ;
        RECT 28.600 166.400 29.000 166.500 ;
        RECT 27.100 166.100 29.000 166.400 ;
        RECT 27.100 166.000 27.500 166.100 ;
        RECT 27.900 165.700 28.300 165.800 ;
        RECT 26.200 165.400 28.300 165.700 ;
        RECT 26.200 161.100 26.600 165.400 ;
        RECT 29.500 165.200 29.800 166.800 ;
        RECT 33.100 166.700 33.500 166.800 ;
        RECT 32.600 166.200 33.000 166.300 ;
        RECT 33.900 166.200 34.300 166.300 ;
        RECT 31.800 165.900 34.300 166.200 ;
        RECT 31.800 165.800 32.200 165.900 ;
        RECT 37.400 165.800 37.800 166.600 ;
        RECT 38.200 165.800 38.600 166.600 ;
        RECT 39.000 166.500 39.700 166.900 ;
        RECT 40.000 166.800 41.800 167.100 ;
        RECT 32.600 165.500 35.400 165.600 ;
        RECT 39.000 165.500 39.300 166.500 ;
        RECT 32.500 165.400 35.400 165.500 ;
        RECT 28.600 164.900 29.800 165.200 ;
        RECT 30.500 165.300 35.400 165.400 ;
        RECT 30.500 165.100 32.900 165.300 ;
        RECT 28.600 164.400 28.900 164.900 ;
        RECT 28.200 164.000 28.900 164.400 ;
        RECT 29.700 164.500 30.100 164.600 ;
        RECT 30.500 164.500 30.800 165.100 ;
        RECT 29.700 164.200 30.800 164.500 ;
        RECT 31.100 164.500 33.800 164.800 ;
        RECT 31.100 164.400 31.500 164.500 ;
        RECT 33.400 164.400 33.800 164.500 ;
        RECT 30.300 163.700 30.700 163.800 ;
        RECT 31.700 163.700 32.100 163.800 ;
        RECT 28.600 163.100 29.000 163.500 ;
        RECT 30.300 163.400 32.100 163.700 ;
        RECT 30.700 163.100 31.000 163.400 ;
        RECT 33.400 163.100 33.800 163.500 ;
        RECT 28.300 161.100 28.900 163.100 ;
        RECT 30.600 161.100 31.000 163.100 ;
        RECT 32.800 162.800 33.800 163.100 ;
        RECT 32.800 161.100 33.200 162.800 ;
        RECT 35.000 161.100 35.400 165.300 ;
        RECT 37.400 165.200 39.300 165.500 ;
        RECT 37.400 163.500 37.700 165.200 ;
        RECT 40.000 164.900 40.300 166.800 ;
        RECT 40.600 166.100 41.000 166.200 ;
        RECT 42.200 166.100 42.600 169.900 ;
        RECT 43.000 167.800 43.400 168.600 ;
        RECT 43.800 167.500 44.200 169.900 ;
        RECT 46.000 169.200 46.400 169.900 ;
        RECT 45.400 168.900 46.400 169.200 ;
        RECT 48.200 168.900 48.600 169.900 ;
        RECT 50.300 169.200 50.900 169.900 ;
        RECT 50.200 168.900 50.900 169.200 ;
        RECT 45.400 168.500 45.800 168.900 ;
        RECT 48.200 168.600 48.500 168.900 ;
        RECT 46.200 168.200 46.600 168.600 ;
        RECT 47.100 168.300 48.500 168.600 ;
        RECT 50.200 168.500 50.600 168.900 ;
        RECT 47.100 168.200 47.500 168.300 ;
        RECT 44.200 167.100 45.000 167.200 ;
        RECT 46.300 167.100 46.600 168.200 ;
        RECT 51.100 167.700 51.500 167.800 ;
        RECT 52.600 167.700 53.000 169.900 ;
        RECT 51.100 167.400 53.000 167.700 ;
        RECT 54.200 167.600 54.600 169.900 ;
        RECT 55.800 167.600 56.200 169.900 ;
        RECT 57.400 167.600 57.800 169.900 ;
        RECT 59.000 167.600 59.400 169.900 ;
        RECT 49.100 167.100 49.500 167.200 ;
        RECT 44.200 166.800 49.700 167.100 ;
        RECT 45.700 166.700 46.100 166.800 ;
        RECT 40.600 165.800 42.600 166.100 ;
        RECT 44.900 166.200 45.300 166.300 ;
        RECT 46.200 166.200 46.600 166.300 ;
        RECT 49.400 166.200 49.700 166.800 ;
        RECT 50.200 166.400 50.600 166.500 ;
        RECT 44.900 165.900 47.400 166.200 ;
        RECT 47.000 165.800 47.400 165.900 ;
        RECT 49.400 165.800 49.800 166.200 ;
        RECT 50.200 166.100 52.100 166.400 ;
        RECT 51.700 166.000 52.100 166.100 ;
        RECT 40.600 165.400 41.000 165.800 ;
        RECT 39.500 164.600 40.300 164.900 ;
        RECT 37.400 161.500 37.800 163.500 ;
        RECT 39.500 161.100 39.900 164.600 ;
        RECT 42.200 161.100 42.600 165.800 ;
        RECT 43.800 165.500 46.600 165.600 ;
        RECT 43.800 165.400 46.700 165.500 ;
        RECT 43.800 165.300 48.700 165.400 ;
        RECT 43.800 161.100 44.200 165.300 ;
        RECT 46.300 165.100 48.700 165.300 ;
        RECT 45.400 164.500 48.100 164.800 ;
        RECT 45.400 164.400 45.800 164.500 ;
        RECT 47.700 164.400 48.100 164.500 ;
        RECT 48.400 164.500 48.700 165.100 ;
        RECT 49.400 165.200 49.700 165.800 ;
        RECT 50.900 165.700 51.300 165.800 ;
        RECT 52.600 165.700 53.000 167.400 ;
        RECT 50.900 165.400 53.000 165.700 ;
        RECT 53.400 167.200 54.600 167.600 ;
        RECT 55.100 167.200 56.200 167.600 ;
        RECT 56.700 167.200 57.800 167.600 ;
        RECT 58.500 167.200 59.400 167.600 ;
        RECT 60.600 167.500 61.000 169.900 ;
        RECT 62.800 169.200 63.200 169.900 ;
        RECT 62.200 168.900 63.200 169.200 ;
        RECT 65.000 168.900 65.400 169.900 ;
        RECT 67.100 169.200 67.700 169.900 ;
        RECT 67.000 168.900 67.700 169.200 ;
        RECT 62.200 168.500 62.600 168.900 ;
        RECT 65.000 168.600 65.300 168.900 ;
        RECT 63.000 168.200 63.400 168.600 ;
        RECT 63.900 168.300 65.300 168.600 ;
        RECT 67.000 168.500 67.400 168.900 ;
        RECT 63.900 168.200 64.300 168.300 ;
        RECT 53.400 165.800 53.800 167.200 ;
        RECT 55.100 166.900 55.500 167.200 ;
        RECT 56.700 166.900 57.100 167.200 ;
        RECT 58.500 166.900 58.900 167.200 ;
        RECT 54.200 166.500 55.500 166.900 ;
        RECT 55.900 166.500 57.100 166.900 ;
        RECT 57.600 166.500 58.900 166.900 ;
        RECT 61.000 167.100 61.800 167.200 ;
        RECT 63.100 167.100 63.400 168.200 ;
        RECT 67.900 167.700 68.300 167.800 ;
        RECT 69.400 167.700 69.800 169.900 ;
        RECT 67.900 167.400 69.800 167.700 ;
        RECT 65.900 167.100 66.300 167.200 ;
        RECT 61.000 166.800 66.500 167.100 ;
        RECT 62.500 166.700 62.900 166.800 ;
        RECT 55.100 165.800 55.500 166.500 ;
        RECT 56.700 165.800 57.100 166.500 ;
        RECT 58.500 165.800 58.900 166.500 ;
        RECT 61.700 166.200 62.100 166.300 ;
        RECT 61.700 165.900 64.200 166.200 ;
        RECT 63.800 165.800 64.200 165.900 ;
        RECT 53.400 165.400 54.600 165.800 ;
        RECT 55.100 165.400 56.200 165.800 ;
        RECT 56.700 165.400 57.800 165.800 ;
        RECT 58.500 165.400 59.400 165.800 ;
        RECT 49.400 164.900 50.600 165.200 ;
        RECT 49.100 164.500 49.500 164.600 ;
        RECT 48.400 164.200 49.500 164.500 ;
        RECT 50.300 164.400 50.600 164.900 ;
        RECT 50.300 164.000 51.000 164.400 ;
        RECT 47.100 163.700 47.500 163.800 ;
        RECT 48.500 163.700 48.900 163.800 ;
        RECT 45.400 163.100 45.800 163.500 ;
        RECT 47.100 163.400 48.900 163.700 ;
        RECT 48.200 163.100 48.500 163.400 ;
        RECT 50.200 163.100 50.600 163.500 ;
        RECT 45.400 162.800 46.400 163.100 ;
        RECT 46.000 161.100 46.400 162.800 ;
        RECT 48.200 161.100 48.600 163.100 ;
        RECT 50.300 161.100 50.900 163.100 ;
        RECT 52.600 161.100 53.000 165.400 ;
        RECT 54.200 161.100 54.600 165.400 ;
        RECT 55.800 161.100 56.200 165.400 ;
        RECT 57.400 161.100 57.800 165.400 ;
        RECT 59.000 161.100 59.400 165.400 ;
        RECT 60.600 165.500 63.400 165.600 ;
        RECT 60.600 165.400 63.500 165.500 ;
        RECT 60.600 165.300 65.500 165.400 ;
        RECT 60.600 161.100 61.000 165.300 ;
        RECT 63.100 165.100 65.500 165.300 ;
        RECT 62.200 164.500 64.900 164.800 ;
        RECT 62.200 164.400 62.600 164.500 ;
        RECT 64.500 164.400 64.900 164.500 ;
        RECT 65.200 164.500 65.500 165.100 ;
        RECT 66.200 165.200 66.500 166.800 ;
        RECT 67.000 166.400 67.400 166.500 ;
        RECT 67.000 166.100 68.900 166.400 ;
        RECT 68.500 166.000 68.900 166.100 ;
        RECT 67.700 165.700 68.100 165.800 ;
        RECT 69.400 165.700 69.800 167.400 ;
        RECT 71.000 167.600 71.400 169.900 ;
        RECT 72.600 167.600 73.000 169.900 ;
        RECT 71.000 167.200 73.000 167.600 ;
        RECT 75.000 167.600 75.400 169.900 ;
        RECT 76.600 167.600 77.000 169.900 ;
        RECT 78.200 167.600 78.600 169.900 ;
        RECT 79.800 167.600 80.200 169.900 ;
        RECT 82.200 167.600 82.600 169.900 ;
        RECT 83.800 167.600 84.200 169.900 ;
        RECT 75.000 167.200 75.900 167.600 ;
        RECT 76.600 167.200 77.700 167.600 ;
        RECT 78.200 167.200 79.300 167.600 ;
        RECT 79.800 167.200 81.000 167.600 ;
        RECT 82.200 167.200 84.200 167.600 ;
        RECT 86.200 167.600 86.600 169.900 ;
        RECT 87.800 167.600 88.200 169.900 ;
        RECT 86.200 167.200 88.200 167.600 ;
        RECT 91.000 167.500 91.400 169.900 ;
        RECT 93.200 169.200 93.600 169.900 ;
        RECT 92.600 168.900 93.600 169.200 ;
        RECT 95.400 168.900 95.800 169.900 ;
        RECT 97.500 169.200 98.100 169.900 ;
        RECT 97.400 168.900 98.100 169.200 ;
        RECT 92.600 168.500 93.000 168.900 ;
        RECT 95.400 168.600 95.700 168.900 ;
        RECT 93.400 168.200 93.800 168.600 ;
        RECT 94.300 168.300 95.700 168.600 ;
        RECT 97.400 168.500 97.800 168.900 ;
        RECT 94.300 168.200 94.700 168.300 ;
        RECT 72.600 165.800 73.000 167.200 ;
        RECT 75.500 166.900 75.900 167.200 ;
        RECT 77.300 166.900 77.700 167.200 ;
        RECT 78.900 166.900 79.300 167.200 ;
        RECT 75.500 166.500 76.800 166.900 ;
        RECT 77.300 166.500 78.500 166.900 ;
        RECT 78.900 166.500 80.200 166.900 ;
        RECT 75.500 165.800 75.900 166.500 ;
        RECT 77.300 165.800 77.700 166.500 ;
        RECT 78.900 165.800 79.300 166.500 ;
        RECT 80.600 165.800 81.000 167.200 ;
        RECT 83.800 165.800 84.200 167.200 ;
        RECT 87.800 166.100 88.200 167.200 ;
        RECT 91.400 167.100 92.200 167.200 ;
        RECT 93.500 167.100 93.800 168.200 ;
        RECT 98.300 167.700 98.700 167.800 ;
        RECT 99.800 167.700 100.200 169.900 ;
        RECT 98.300 167.400 100.200 167.700 ;
        RECT 96.300 167.100 96.700 167.200 ;
        RECT 91.400 166.800 96.900 167.100 ;
        RECT 92.900 166.700 93.300 166.800 ;
        RECT 92.100 166.200 92.500 166.300 ;
        RECT 88.600 166.100 89.000 166.200 ;
        RECT 87.800 165.800 89.000 166.100 ;
        RECT 92.100 165.900 94.600 166.200 ;
        RECT 94.200 165.800 94.600 165.900 ;
        RECT 67.700 165.400 69.800 165.700 ;
        RECT 66.200 164.900 67.400 165.200 ;
        RECT 65.900 164.500 66.300 164.600 ;
        RECT 65.200 164.200 66.300 164.500 ;
        RECT 67.100 164.400 67.400 164.900 ;
        RECT 67.100 164.200 67.800 164.400 ;
        RECT 67.100 164.000 68.200 164.200 ;
        RECT 67.500 163.800 68.200 164.000 ;
        RECT 63.900 163.700 64.300 163.800 ;
        RECT 65.300 163.700 65.700 163.800 ;
        RECT 62.200 163.100 62.600 163.500 ;
        RECT 63.900 163.400 65.700 163.700 ;
        RECT 65.000 163.100 65.300 163.400 ;
        RECT 67.000 163.100 67.400 163.500 ;
        RECT 62.200 162.800 63.200 163.100 ;
        RECT 62.800 161.100 63.200 162.800 ;
        RECT 65.000 161.100 65.400 163.100 ;
        RECT 67.100 161.100 67.700 163.100 ;
        RECT 69.400 161.100 69.800 165.400 ;
        RECT 71.000 165.400 73.000 165.800 ;
        RECT 71.000 161.100 71.400 165.400 ;
        RECT 72.600 161.100 73.000 165.400 ;
        RECT 75.000 165.400 75.900 165.800 ;
        RECT 76.600 165.400 77.700 165.800 ;
        RECT 78.200 165.400 79.300 165.800 ;
        RECT 79.800 165.400 81.000 165.800 ;
        RECT 82.200 165.400 84.200 165.800 ;
        RECT 75.000 161.100 75.400 165.400 ;
        RECT 76.600 161.100 77.000 165.400 ;
        RECT 78.200 161.100 78.600 165.400 ;
        RECT 79.800 161.100 80.200 165.400 ;
        RECT 82.200 161.100 82.600 165.400 ;
        RECT 83.800 161.100 84.200 165.400 ;
        RECT 86.200 165.400 88.200 165.800 ;
        RECT 86.200 161.100 86.600 165.400 ;
        RECT 87.800 161.100 88.200 165.400 ;
        RECT 91.000 165.500 93.800 165.600 ;
        RECT 91.000 165.400 93.900 165.500 ;
        RECT 91.000 165.300 95.900 165.400 ;
        RECT 91.000 161.100 91.400 165.300 ;
        RECT 93.500 165.100 95.900 165.300 ;
        RECT 92.600 164.500 95.300 164.800 ;
        RECT 92.600 164.400 93.000 164.500 ;
        RECT 94.900 164.400 95.300 164.500 ;
        RECT 95.600 164.500 95.900 165.100 ;
        RECT 96.600 165.200 96.900 166.800 ;
        RECT 97.400 166.400 97.800 166.500 ;
        RECT 97.400 166.100 99.300 166.400 ;
        RECT 98.900 166.000 99.300 166.100 ;
        RECT 98.100 165.700 98.500 165.800 ;
        RECT 99.800 165.700 100.200 167.400 ;
        RECT 100.600 168.500 101.000 169.500 ;
        RECT 100.600 167.400 100.900 168.500 ;
        RECT 102.700 168.000 103.100 169.500 ;
        RECT 102.700 167.700 103.500 168.000 ;
        RECT 103.100 167.500 103.500 167.700 ;
        RECT 100.600 167.100 102.700 167.400 ;
        RECT 102.200 166.900 102.700 167.100 ;
        RECT 103.200 167.200 103.500 167.500 ;
        RECT 103.200 167.100 104.200 167.200 ;
        RECT 104.600 167.100 105.000 167.200 ;
        RECT 100.600 165.800 101.000 166.600 ;
        RECT 101.400 165.800 101.800 166.600 ;
        RECT 102.200 166.500 102.900 166.900 ;
        RECT 103.200 166.800 105.000 167.100 ;
        RECT 98.100 165.400 100.200 165.700 ;
        RECT 102.200 165.500 102.500 166.500 ;
        RECT 96.600 164.900 97.800 165.200 ;
        RECT 96.300 164.500 96.700 164.600 ;
        RECT 95.600 164.200 96.700 164.500 ;
        RECT 97.500 164.400 97.800 164.900 ;
        RECT 97.500 164.000 98.200 164.400 ;
        RECT 94.300 163.700 94.700 163.800 ;
        RECT 95.700 163.700 96.100 163.800 ;
        RECT 92.600 163.100 93.000 163.500 ;
        RECT 94.300 163.400 96.100 163.700 ;
        RECT 95.400 163.100 95.700 163.400 ;
        RECT 97.400 163.100 97.800 163.500 ;
        RECT 92.600 162.800 93.600 163.100 ;
        RECT 93.200 161.100 93.600 162.800 ;
        RECT 95.400 161.100 95.800 163.100 ;
        RECT 97.500 161.100 98.100 163.100 ;
        RECT 99.800 161.100 100.200 165.400 ;
        RECT 100.600 165.200 102.500 165.500 ;
        RECT 100.600 163.500 100.900 165.200 ;
        RECT 103.200 164.900 103.500 166.800 ;
        RECT 103.800 166.100 104.200 166.200 ;
        RECT 105.400 166.100 105.800 169.900 ;
        RECT 106.200 168.100 106.600 168.600 ;
        RECT 107.000 168.100 107.400 169.900 ;
        RECT 109.100 169.200 109.700 169.900 ;
        RECT 109.100 168.900 109.800 169.200 ;
        RECT 111.400 168.900 111.800 169.900 ;
        RECT 113.600 169.200 114.000 169.900 ;
        RECT 113.600 168.900 114.600 169.200 ;
        RECT 109.400 168.500 109.800 168.900 ;
        RECT 111.500 168.600 111.800 168.900 ;
        RECT 111.500 168.300 112.900 168.600 ;
        RECT 112.500 168.200 112.900 168.300 ;
        RECT 113.400 168.200 113.800 168.600 ;
        RECT 114.200 168.500 114.600 168.900 ;
        RECT 106.200 167.800 107.400 168.100 ;
        RECT 103.800 165.800 105.800 166.100 ;
        RECT 103.800 165.400 104.200 165.800 ;
        RECT 102.700 164.600 103.500 164.900 ;
        RECT 100.600 161.500 101.000 163.500 ;
        RECT 102.700 161.100 103.100 164.600 ;
        RECT 105.400 161.100 105.800 165.800 ;
        RECT 107.000 167.700 107.400 167.800 ;
        RECT 108.500 167.700 108.900 167.800 ;
        RECT 107.000 167.400 108.900 167.700 ;
        RECT 107.000 165.700 107.400 167.400 ;
        RECT 110.500 167.100 110.900 167.200 ;
        RECT 112.600 167.100 113.000 167.200 ;
        RECT 113.400 167.100 113.700 168.200 ;
        RECT 115.800 167.500 116.200 169.900 ;
        RECT 117.400 168.000 117.800 169.900 ;
        RECT 117.300 167.600 117.800 168.000 ;
        RECT 115.000 167.100 115.800 167.200 ;
        RECT 110.300 166.800 115.800 167.100 ;
        RECT 109.400 166.400 109.800 166.500 ;
        RECT 107.900 166.100 109.800 166.400 ;
        RECT 107.900 166.000 108.300 166.100 ;
        RECT 108.700 165.700 109.100 165.800 ;
        RECT 107.000 165.400 109.100 165.700 ;
        RECT 107.000 161.100 107.400 165.400 ;
        RECT 110.300 165.200 110.600 166.800 ;
        RECT 113.900 166.700 114.300 166.800 ;
        RECT 114.700 166.200 115.100 166.300 ;
        RECT 111.800 166.100 112.200 166.200 ;
        RECT 112.600 166.100 115.100 166.200 ;
        RECT 111.800 165.900 115.100 166.100 ;
        RECT 111.800 165.800 113.000 165.900 ;
        RECT 113.400 165.500 116.200 165.600 ;
        RECT 113.300 165.400 116.200 165.500 ;
        RECT 109.400 164.900 110.600 165.200 ;
        RECT 111.300 165.300 116.200 165.400 ;
        RECT 111.300 165.100 113.700 165.300 ;
        RECT 109.400 164.400 109.700 164.900 ;
        RECT 109.000 164.000 109.700 164.400 ;
        RECT 110.500 164.500 110.900 164.600 ;
        RECT 111.300 164.500 111.600 165.100 ;
        RECT 110.500 164.200 111.600 164.500 ;
        RECT 111.900 164.500 114.600 164.800 ;
        RECT 111.900 164.400 112.300 164.500 ;
        RECT 114.200 164.400 114.600 164.500 ;
        RECT 111.100 163.700 111.500 163.800 ;
        RECT 112.500 163.700 112.900 163.800 ;
        RECT 109.400 163.100 109.800 163.500 ;
        RECT 111.100 163.400 112.900 163.700 ;
        RECT 111.500 163.100 111.800 163.400 ;
        RECT 114.200 163.100 114.600 163.500 ;
        RECT 109.100 161.100 109.700 163.100 ;
        RECT 111.400 161.100 111.800 163.100 ;
        RECT 113.600 162.800 114.600 163.100 ;
        RECT 113.600 161.100 114.000 162.800 ;
        RECT 115.800 161.100 116.200 165.300 ;
        RECT 117.300 165.400 117.700 167.600 ;
        RECT 118.200 167.300 118.600 169.900 ;
        RECT 121.400 168.300 121.800 169.900 ;
        RECT 122.200 168.500 122.600 169.900 ;
        RECT 123.000 168.500 123.400 169.900 ;
        RECT 123.800 168.500 124.200 169.900 ;
        RECT 124.600 168.500 125.000 169.900 ;
        RECT 126.200 168.500 126.600 169.900 ;
        RECT 127.800 168.500 128.200 169.900 ;
        RECT 128.600 168.500 129.000 169.900 ;
        RECT 129.400 168.500 129.800 169.900 ;
        RECT 120.600 167.900 121.800 168.300 ;
        RECT 130.200 168.300 130.600 169.900 ;
        RECT 120.600 167.600 121.000 167.900 ;
        RECT 118.000 167.000 118.600 167.300 ;
        RECT 120.100 167.300 121.000 167.600 ;
        RECT 123.000 167.800 123.500 168.200 ;
        RECT 125.000 167.800 125.800 168.200 ;
        RECT 126.200 167.900 128.500 168.200 ;
        RECT 130.200 167.900 131.500 168.300 ;
        RECT 126.200 167.800 126.600 167.900 ;
        RECT 118.000 166.000 118.300 167.000 ;
        RECT 120.100 166.700 120.500 167.300 ;
        RECT 118.600 166.300 120.500 166.700 ;
        RECT 123.000 166.400 123.400 167.800 ;
        RECT 126.200 167.400 126.600 167.500 ;
        RECT 124.400 167.100 126.600 167.400 ;
        RECT 124.400 167.000 124.800 167.100 ;
        RECT 127.000 166.800 127.400 167.600 ;
        RECT 128.100 166.700 128.500 167.900 ;
        RECT 131.100 167.600 131.500 167.900 ;
        RECT 131.100 167.200 132.600 167.600 ;
        RECT 133.400 166.900 133.800 169.900 ;
        RECT 124.600 166.300 126.200 166.700 ;
        RECT 128.100 166.300 129.100 166.700 ;
        RECT 129.400 166.500 133.800 166.900 ;
        RECT 118.000 165.700 118.400 166.000 ;
        RECT 117.300 165.000 117.800 165.400 ;
        RECT 117.400 161.100 117.800 165.000 ;
        RECT 118.100 164.800 118.400 165.700 ;
        RECT 118.100 164.500 122.600 164.800 ;
        RECT 118.100 163.700 118.400 164.500 ;
        RECT 122.200 164.400 122.600 164.500 ;
        RECT 123.800 164.500 128.100 164.800 ;
        RECT 123.800 164.400 124.200 164.500 ;
        RECT 119.700 163.800 121.000 164.200 ;
        RECT 118.100 163.400 119.400 163.700 ;
        RECT 119.000 161.100 119.400 163.400 ;
        RECT 120.600 161.100 121.000 163.800 ;
        RECT 121.300 163.400 123.400 163.800 ;
        RECT 122.200 161.100 122.600 162.500 ;
        RECT 123.000 161.100 123.400 162.500 ;
        RECT 123.800 161.100 124.200 162.500 ;
        RECT 124.600 161.100 125.000 164.200 ;
        RECT 126.200 163.800 127.500 164.200 ;
        RECT 127.800 164.100 128.100 164.500 ;
        RECT 128.600 164.700 129.000 164.800 ;
        RECT 128.600 164.500 131.300 164.700 ;
        RECT 128.600 164.400 131.700 164.500 ;
        RECT 131.000 164.100 131.700 164.400 ;
        RECT 127.800 163.800 130.700 164.100 ;
        RECT 132.200 164.000 133.000 164.400 ;
        RECT 132.200 163.800 132.500 164.000 ;
        RECT 126.200 161.100 126.600 163.500 ;
        RECT 127.800 161.100 128.200 163.500 ;
        RECT 130.400 163.400 132.500 163.800 ;
        RECT 133.400 163.700 133.800 166.500 ;
        RECT 132.800 163.400 133.800 163.700 ;
        RECT 135.800 166.900 136.200 169.900 ;
        RECT 139.000 168.300 139.400 169.900 ;
        RECT 139.800 168.500 140.200 169.900 ;
        RECT 140.600 168.500 141.000 169.900 ;
        RECT 141.400 168.500 141.800 169.900 ;
        RECT 143.000 168.500 143.400 169.900 ;
        RECT 144.600 168.500 145.000 169.900 ;
        RECT 145.400 168.500 145.800 169.900 ;
        RECT 146.200 168.500 146.600 169.900 ;
        RECT 147.000 168.500 147.400 169.900 ;
        RECT 138.100 167.900 139.400 168.300 ;
        RECT 147.800 168.300 148.200 169.900 ;
        RECT 141.100 167.900 143.400 168.200 ;
        RECT 138.100 167.600 138.500 167.900 ;
        RECT 137.000 167.200 138.500 167.600 ;
        RECT 135.800 166.500 140.200 166.900 ;
        RECT 141.100 166.700 141.500 167.900 ;
        RECT 143.000 167.800 143.400 167.900 ;
        RECT 143.800 167.800 144.600 168.200 ;
        RECT 146.100 167.800 146.600 168.200 ;
        RECT 147.800 167.900 149.000 168.300 ;
        RECT 142.200 166.800 142.600 167.600 ;
        RECT 143.000 167.400 143.400 167.500 ;
        RECT 143.000 167.100 145.200 167.400 ;
        RECT 144.800 167.000 145.200 167.100 ;
        RECT 135.800 163.700 136.200 166.500 ;
        RECT 140.500 166.300 141.500 166.700 ;
        RECT 143.400 166.300 145.000 166.700 ;
        RECT 146.200 166.400 146.600 167.800 ;
        RECT 148.600 167.600 149.000 167.900 ;
        RECT 148.600 167.300 149.500 167.600 ;
        RECT 149.100 166.700 149.500 167.300 ;
        RECT 151.000 167.300 151.400 169.900 ;
        RECT 151.800 168.000 152.200 169.900 ;
        RECT 151.800 167.600 152.300 168.000 ;
        RECT 151.000 167.000 151.600 167.300 ;
        RECT 149.100 166.300 151.000 166.700 ;
        RECT 151.300 166.000 151.600 167.000 ;
        RECT 151.200 165.700 151.600 166.000 ;
        RECT 151.900 166.100 152.300 167.600 ;
        RECT 153.400 167.600 153.800 169.900 ;
        RECT 153.400 167.300 154.500 167.600 ;
        RECT 155.800 167.500 156.200 169.900 ;
        RECT 158.000 169.200 158.400 169.900 ;
        RECT 157.400 168.900 158.400 169.200 ;
        RECT 160.200 168.900 160.600 169.900 ;
        RECT 162.300 169.200 162.900 169.900 ;
        RECT 162.200 168.900 162.900 169.200 ;
        RECT 157.400 168.500 157.800 168.900 ;
        RECT 160.200 168.600 160.500 168.900 ;
        RECT 158.200 168.200 158.600 168.600 ;
        RECT 159.100 168.300 160.500 168.600 ;
        RECT 162.200 168.500 162.600 168.900 ;
        RECT 159.100 168.200 159.500 168.300 ;
        RECT 153.400 166.100 153.800 166.600 ;
        RECT 151.900 165.800 153.800 166.100 ;
        RECT 154.200 165.800 154.500 167.300 ;
        RECT 156.200 167.100 157.000 167.200 ;
        RECT 158.300 167.100 158.600 168.200 ;
        RECT 163.100 167.700 163.500 167.800 ;
        RECT 164.600 167.700 165.000 169.900 ;
        RECT 163.100 167.400 165.000 167.700 ;
        RECT 161.100 167.100 161.500 167.200 ;
        RECT 156.200 166.800 161.700 167.100 ;
        RECT 157.700 166.700 158.100 166.800 ;
        RECT 156.900 166.200 157.300 166.300 ;
        RECT 156.900 165.900 159.400 166.200 ;
        RECT 159.000 165.800 159.400 165.900 ;
        RECT 151.200 164.800 151.500 165.700 ;
        RECT 151.900 165.400 152.300 165.800 ;
        RECT 140.600 164.700 141.000 164.800 ;
        RECT 138.300 164.500 141.000 164.700 ;
        RECT 137.900 164.400 141.000 164.500 ;
        RECT 141.500 164.500 145.800 164.800 ;
        RECT 136.600 164.000 137.400 164.400 ;
        RECT 137.900 164.100 138.600 164.400 ;
        RECT 141.500 164.100 141.800 164.500 ;
        RECT 145.400 164.400 145.800 164.500 ;
        RECT 147.000 164.500 151.500 164.800 ;
        RECT 147.000 164.400 147.400 164.500 ;
        RECT 137.100 163.800 137.400 164.000 ;
        RECT 138.900 163.800 141.800 164.100 ;
        RECT 142.100 163.800 143.400 164.200 ;
        RECT 135.800 163.400 136.800 163.700 ;
        RECT 137.100 163.400 139.200 163.800 ;
        RECT 128.600 161.100 129.000 162.500 ;
        RECT 129.400 161.100 129.800 162.500 ;
        RECT 131.000 161.100 131.400 163.400 ;
        RECT 132.800 163.100 133.100 163.400 ;
        RECT 132.600 162.800 133.100 163.100 ;
        RECT 136.500 163.100 136.800 163.400 ;
        RECT 136.500 162.800 137.000 163.100 ;
        RECT 132.600 161.100 133.000 162.800 ;
        RECT 136.600 161.100 137.000 162.800 ;
        RECT 138.200 161.100 138.600 163.400 ;
        RECT 139.800 161.100 140.200 162.500 ;
        RECT 140.600 161.100 141.000 162.500 ;
        RECT 141.400 161.100 141.800 163.500 ;
        RECT 143.000 161.100 143.400 163.500 ;
        RECT 144.600 161.100 145.000 164.200 ;
        RECT 148.600 163.800 149.900 164.200 ;
        RECT 146.200 163.400 148.300 163.800 ;
        RECT 145.400 161.100 145.800 162.500 ;
        RECT 146.200 161.100 146.600 162.500 ;
        RECT 147.000 161.100 147.400 162.500 ;
        RECT 148.600 161.100 149.000 163.800 ;
        RECT 151.200 163.700 151.500 164.500 ;
        RECT 150.200 163.400 151.500 163.700 ;
        RECT 151.800 165.000 152.300 165.400 ;
        RECT 154.200 165.400 154.800 165.800 ;
        RECT 155.800 165.500 158.600 165.600 ;
        RECT 155.800 165.400 158.700 165.500 ;
        RECT 154.200 165.100 154.500 165.400 ;
        RECT 150.200 161.100 150.600 163.400 ;
        RECT 151.800 161.100 152.200 165.000 ;
        RECT 153.400 164.800 154.500 165.100 ;
        RECT 155.800 165.300 160.700 165.400 ;
        RECT 153.400 161.100 153.800 164.800 ;
        RECT 155.800 161.100 156.200 165.300 ;
        RECT 158.300 165.100 160.700 165.300 ;
        RECT 157.400 164.500 160.100 164.800 ;
        RECT 157.400 164.400 157.800 164.500 ;
        RECT 159.700 164.400 160.100 164.500 ;
        RECT 160.400 164.500 160.700 165.100 ;
        RECT 161.400 165.200 161.700 166.800 ;
        RECT 162.200 166.400 162.600 166.500 ;
        RECT 162.200 166.100 164.100 166.400 ;
        RECT 163.700 166.000 164.100 166.100 ;
        RECT 162.900 165.700 163.300 165.800 ;
        RECT 164.600 165.700 165.000 167.400 ;
        RECT 165.400 168.500 165.800 169.500 ;
        RECT 165.400 167.400 165.700 168.500 ;
        RECT 167.500 168.000 167.900 169.500 ;
        RECT 170.200 168.500 170.600 169.500 ;
        RECT 167.500 167.700 168.300 168.000 ;
        RECT 167.900 167.500 168.300 167.700 ;
        RECT 165.400 167.100 167.500 167.400 ;
        RECT 167.000 166.900 167.500 167.100 ;
        RECT 168.000 167.200 168.300 167.500 ;
        RECT 170.200 167.400 170.500 168.500 ;
        RECT 172.300 168.000 172.700 169.500 ;
        RECT 172.300 167.700 173.100 168.000 ;
        RECT 172.700 167.500 173.100 167.700 ;
        RECT 165.400 165.800 165.800 166.600 ;
        RECT 166.200 165.800 166.600 166.600 ;
        RECT 167.000 166.500 167.700 166.900 ;
        RECT 168.000 166.800 169.000 167.200 ;
        RECT 170.200 167.100 172.300 167.400 ;
        RECT 171.800 166.900 172.300 167.100 ;
        RECT 172.800 167.200 173.100 167.500 ;
        RECT 175.000 167.600 175.400 169.900 ;
        RECT 177.400 167.600 177.800 169.900 ;
        RECT 175.000 167.300 176.100 167.600 ;
        RECT 177.400 167.300 178.500 167.600 ;
        RECT 162.900 165.400 165.000 165.700 ;
        RECT 167.000 165.500 167.300 166.500 ;
        RECT 161.400 164.900 162.600 165.200 ;
        RECT 161.100 164.500 161.500 164.600 ;
        RECT 160.400 164.200 161.500 164.500 ;
        RECT 162.300 164.400 162.600 164.900 ;
        RECT 162.300 164.000 163.000 164.400 ;
        RECT 159.100 163.700 159.500 163.800 ;
        RECT 160.500 163.700 160.900 163.800 ;
        RECT 157.400 163.100 157.800 163.500 ;
        RECT 159.100 163.400 160.900 163.700 ;
        RECT 160.200 163.100 160.500 163.400 ;
        RECT 162.200 163.100 162.600 163.500 ;
        RECT 157.400 162.800 158.400 163.100 ;
        RECT 158.000 161.100 158.400 162.800 ;
        RECT 160.200 161.100 160.600 163.100 ;
        RECT 162.300 161.100 162.900 163.100 ;
        RECT 164.600 161.100 165.000 165.400 ;
        RECT 165.400 165.200 167.300 165.500 ;
        RECT 165.400 163.500 165.700 165.200 ;
        RECT 168.000 164.900 168.300 166.800 ;
        RECT 168.600 165.400 169.000 166.200 ;
        RECT 170.200 165.800 170.600 166.600 ;
        RECT 171.000 165.800 171.400 166.600 ;
        RECT 171.800 166.500 172.500 166.900 ;
        RECT 172.800 166.800 173.800 167.200 ;
        RECT 171.800 165.500 172.100 166.500 ;
        RECT 167.500 164.600 168.300 164.900 ;
        RECT 170.200 165.200 172.100 165.500 ;
        RECT 165.400 161.500 165.800 163.500 ;
        RECT 167.500 162.200 167.900 164.600 ;
        RECT 170.200 163.500 170.500 165.200 ;
        RECT 172.800 164.900 173.100 166.800 ;
        RECT 173.400 165.400 173.800 166.200 ;
        RECT 174.200 166.100 174.600 166.200 ;
        RECT 175.000 166.100 175.400 166.600 ;
        RECT 174.200 165.800 175.400 166.100 ;
        RECT 175.800 165.800 176.100 167.300 ;
        RECT 177.400 165.800 177.800 166.600 ;
        RECT 178.200 165.800 178.500 167.300 ;
        RECT 175.800 165.400 176.400 165.800 ;
        RECT 178.200 165.400 178.800 165.800 ;
        RECT 175.800 165.100 176.100 165.400 ;
        RECT 178.200 165.100 178.500 165.400 ;
        RECT 172.300 164.600 173.100 164.900 ;
        RECT 175.000 164.800 176.100 165.100 ;
        RECT 177.400 164.800 178.500 165.100 ;
        RECT 167.500 161.800 168.200 162.200 ;
        RECT 167.500 161.100 167.900 161.800 ;
        RECT 170.200 161.500 170.600 163.500 ;
        RECT 172.300 162.200 172.700 164.600 ;
        RECT 172.300 161.800 173.000 162.200 ;
        RECT 172.300 161.100 172.700 161.800 ;
        RECT 175.000 161.100 175.400 164.800 ;
        RECT 177.400 161.100 177.800 164.800 ;
        RECT 0.600 155.700 1.000 159.900 ;
        RECT 2.800 158.200 3.200 159.900 ;
        RECT 2.200 157.900 3.200 158.200 ;
        RECT 5.000 157.900 5.400 159.900 ;
        RECT 7.100 157.900 7.700 159.900 ;
        RECT 2.200 157.500 2.600 157.900 ;
        RECT 5.000 157.600 5.300 157.900 ;
        RECT 3.900 157.300 5.700 157.600 ;
        RECT 7.000 157.500 7.400 157.900 ;
        RECT 3.900 157.200 4.300 157.300 ;
        RECT 5.300 157.200 5.700 157.300 ;
        RECT 9.400 157.100 9.800 159.900 ;
        RECT 10.200 157.100 10.600 157.200 ;
        RECT 2.200 156.500 2.600 156.600 ;
        RECT 4.500 156.500 4.900 156.600 ;
        RECT 2.200 156.200 4.900 156.500 ;
        RECT 5.200 156.500 6.300 156.800 ;
        RECT 5.200 155.900 5.500 156.500 ;
        RECT 5.900 156.400 6.300 156.500 ;
        RECT 7.100 156.600 7.800 157.000 ;
        RECT 9.400 156.800 10.600 157.100 ;
        RECT 7.100 156.100 7.400 156.600 ;
        RECT 3.100 155.700 5.500 155.900 ;
        RECT 0.600 155.600 5.500 155.700 ;
        RECT 6.200 155.800 7.400 156.100 ;
        RECT 0.600 155.500 3.500 155.600 ;
        RECT 0.600 155.400 3.400 155.500 ;
        RECT 6.200 155.200 6.500 155.800 ;
        RECT 9.400 155.600 9.800 156.800 ;
        RECT 7.700 155.300 9.800 155.600 ;
        RECT 7.700 155.200 8.100 155.300 ;
        RECT 3.800 155.100 4.200 155.200 ;
        RECT 1.700 154.800 4.200 155.100 ;
        RECT 6.200 154.800 6.600 155.200 ;
        RECT 8.500 154.900 8.900 155.000 ;
        RECT 1.700 154.700 2.100 154.800 ;
        RECT 2.500 154.200 2.900 154.300 ;
        RECT 6.200 154.200 6.500 154.800 ;
        RECT 7.000 154.600 8.900 154.900 ;
        RECT 7.000 154.500 7.400 154.600 ;
        RECT 1.000 153.900 6.500 154.200 ;
        RECT 1.000 153.800 1.800 153.900 ;
        RECT 0.600 151.100 1.000 153.500 ;
        RECT 3.100 152.800 3.400 153.900 ;
        RECT 5.900 153.800 6.300 153.900 ;
        RECT 9.400 153.600 9.800 155.300 ;
        RECT 7.900 153.300 9.800 153.600 ;
        RECT 7.900 153.200 8.300 153.300 ;
        RECT 2.200 152.100 2.600 152.500 ;
        RECT 3.000 152.400 3.400 152.800 ;
        RECT 3.900 152.700 4.300 152.800 ;
        RECT 3.900 152.400 5.300 152.700 ;
        RECT 5.000 152.100 5.300 152.400 ;
        RECT 7.000 152.100 7.400 152.500 ;
        RECT 2.200 151.800 3.200 152.100 ;
        RECT 2.800 151.100 3.200 151.800 ;
        RECT 5.000 151.100 5.400 152.100 ;
        RECT 7.000 151.800 7.700 152.100 ;
        RECT 7.100 151.100 7.700 151.800 ;
        RECT 9.400 151.100 9.800 153.300 ;
        RECT 11.000 155.100 11.400 159.900 ;
        RECT 13.700 156.400 14.100 159.900 ;
        RECT 15.800 157.500 16.200 159.500 ;
        RECT 13.300 156.100 14.100 156.400 ;
        RECT 12.600 155.100 13.000 155.600 ;
        RECT 11.000 154.800 13.000 155.100 ;
        RECT 10.200 152.400 10.600 153.200 ;
        RECT 11.000 151.100 11.400 154.800 ;
        RECT 13.300 154.200 13.600 156.100 ;
        RECT 15.900 155.800 16.200 157.500 ;
        RECT 14.300 155.500 16.200 155.800 ;
        RECT 14.300 154.500 14.600 155.500 ;
        RECT 11.800 154.100 12.200 154.200 ;
        RECT 12.600 154.100 13.600 154.200 ;
        RECT 13.900 154.100 14.600 154.500 ;
        RECT 15.000 154.400 15.400 155.200 ;
        RECT 15.800 154.400 16.200 155.200 ;
        RECT 11.800 153.800 13.600 154.100 ;
        RECT 13.300 153.500 13.600 153.800 ;
        RECT 14.100 153.900 14.600 154.100 ;
        RECT 14.100 153.600 16.200 153.900 ;
        RECT 13.300 153.300 13.700 153.500 ;
        RECT 13.300 153.000 14.100 153.300 ;
        RECT 13.700 151.500 14.100 153.000 ;
        RECT 15.900 152.500 16.200 153.600 ;
        RECT 16.600 153.400 17.000 154.200 ;
        RECT 17.400 153.100 17.800 159.900 ;
        RECT 19.000 157.500 19.400 159.500 ;
        RECT 21.100 159.200 21.500 159.900 ;
        RECT 20.600 158.800 21.500 159.200 ;
        RECT 18.200 155.800 18.600 156.600 ;
        RECT 19.000 155.800 19.300 157.500 ;
        RECT 21.100 156.400 21.500 158.800 ;
        RECT 21.100 156.100 21.900 156.400 ;
        RECT 19.000 155.500 20.900 155.800 ;
        RECT 19.000 154.400 19.400 155.200 ;
        RECT 19.800 154.400 20.200 155.200 ;
        RECT 20.600 154.500 20.900 155.500 ;
        RECT 20.600 154.100 21.300 154.500 ;
        RECT 21.600 154.200 21.900 156.100 ;
        RECT 22.200 155.100 22.600 155.600 ;
        RECT 23.800 155.100 24.200 159.900 ;
        RECT 22.200 154.800 24.200 155.100 ;
        RECT 20.600 153.900 21.100 154.100 ;
        RECT 19.000 153.600 21.100 153.900 ;
        RECT 21.600 153.800 22.600 154.200 ;
        RECT 17.400 152.800 18.300 153.100 ;
        RECT 15.800 151.500 16.200 152.500 ;
        RECT 17.900 152.200 18.300 152.800 ;
        RECT 19.000 152.500 19.300 153.600 ;
        RECT 21.600 153.500 21.900 153.800 ;
        RECT 21.500 153.300 21.900 153.500 ;
        RECT 21.100 153.000 21.900 153.300 ;
        RECT 17.900 151.800 18.600 152.200 ;
        RECT 17.900 151.100 18.300 151.800 ;
        RECT 19.000 151.500 19.400 152.500 ;
        RECT 21.100 151.500 21.500 153.000 ;
        RECT 23.800 151.100 24.200 154.800 ;
        RECT 25.400 154.100 25.800 154.200 ;
        RECT 24.600 153.800 25.800 154.100 ;
        RECT 24.600 153.200 24.900 153.800 ;
        RECT 25.400 153.400 25.800 153.800 ;
        RECT 24.600 152.400 25.000 153.200 ;
        RECT 26.200 153.100 26.600 159.900 ;
        RECT 27.000 155.800 27.400 156.600 ;
        RECT 28.600 155.600 29.000 159.900 ;
        RECT 30.200 155.600 30.600 159.900 ;
        RECT 31.800 155.600 32.200 159.900 ;
        RECT 33.400 155.600 33.800 159.900 ;
        RECT 27.800 155.200 29.000 155.600 ;
        RECT 29.500 155.200 30.600 155.600 ;
        RECT 31.100 155.200 32.200 155.600 ;
        RECT 32.900 155.200 33.800 155.600 ;
        RECT 36.600 155.700 37.000 159.900 ;
        RECT 38.800 158.200 39.200 159.900 ;
        RECT 38.200 157.900 39.200 158.200 ;
        RECT 41.000 157.900 41.400 159.900 ;
        RECT 43.100 157.900 43.700 159.900 ;
        RECT 38.200 157.500 38.600 157.900 ;
        RECT 41.000 157.600 41.300 157.900 ;
        RECT 39.900 157.300 41.700 157.600 ;
        RECT 43.000 157.500 43.400 157.900 ;
        RECT 39.900 157.200 40.300 157.300 ;
        RECT 41.300 157.200 41.700 157.300 ;
        RECT 38.200 156.500 38.600 156.600 ;
        RECT 40.500 156.500 40.900 156.600 ;
        RECT 38.200 156.200 40.900 156.500 ;
        RECT 41.200 156.500 42.300 156.800 ;
        RECT 41.200 155.900 41.500 156.500 ;
        RECT 41.900 156.400 42.300 156.500 ;
        RECT 43.100 156.600 43.800 157.000 ;
        RECT 43.100 156.100 43.400 156.600 ;
        RECT 39.100 155.700 41.500 155.900 ;
        RECT 36.600 155.600 41.500 155.700 ;
        RECT 42.200 155.800 43.400 156.100 ;
        RECT 36.600 155.500 39.500 155.600 ;
        RECT 36.600 155.400 39.400 155.500 ;
        RECT 42.200 155.200 42.500 155.800 ;
        RECT 45.400 155.600 45.800 159.900 ;
        RECT 47.500 156.300 47.900 159.900 ;
        RECT 47.000 155.900 47.900 156.300 ;
        RECT 48.600 155.900 49.000 159.900 ;
        RECT 49.400 156.200 49.800 159.900 ;
        RECT 51.000 156.200 51.400 159.900 ;
        RECT 49.400 155.900 51.400 156.200 ;
        RECT 51.800 157.500 52.200 159.500 ;
        RECT 53.900 158.200 54.300 159.900 ;
        RECT 53.400 157.800 54.300 158.200 ;
        RECT 43.700 155.300 45.800 155.600 ;
        RECT 43.700 155.200 44.100 155.300 ;
        RECT 27.800 153.800 28.200 155.200 ;
        RECT 29.500 154.500 29.900 155.200 ;
        RECT 31.100 154.500 31.500 155.200 ;
        RECT 32.900 154.500 33.300 155.200 ;
        RECT 39.800 155.100 40.200 155.200 ;
        RECT 37.700 154.800 40.200 155.100 ;
        RECT 42.200 154.800 42.600 155.200 ;
        RECT 44.500 154.900 44.900 155.000 ;
        RECT 37.700 154.700 38.100 154.800 ;
        RECT 28.600 154.100 29.900 154.500 ;
        RECT 30.300 154.100 31.500 154.500 ;
        RECT 32.000 154.100 33.300 154.500 ;
        RECT 38.500 154.200 38.900 154.300 ;
        RECT 42.200 154.200 42.500 154.800 ;
        RECT 43.000 154.600 44.900 154.900 ;
        RECT 43.000 154.500 43.400 154.600 ;
        RECT 29.500 153.800 29.900 154.100 ;
        RECT 31.100 153.800 31.500 154.100 ;
        RECT 32.900 153.800 33.300 154.100 ;
        RECT 35.800 154.100 36.200 154.200 ;
        RECT 37.000 154.100 42.500 154.200 ;
        RECT 35.800 153.900 42.500 154.100 ;
        RECT 35.800 153.800 37.800 153.900 ;
        RECT 27.800 153.400 29.000 153.800 ;
        RECT 29.500 153.400 30.600 153.800 ;
        RECT 31.100 153.400 32.200 153.800 ;
        RECT 32.900 153.400 33.800 153.800 ;
        RECT 26.200 152.800 27.100 153.100 ;
        RECT 26.700 152.200 27.100 152.800 ;
        RECT 26.700 151.800 27.400 152.200 ;
        RECT 26.700 151.100 27.100 151.800 ;
        RECT 28.600 151.100 29.000 153.400 ;
        RECT 30.200 151.100 30.600 153.400 ;
        RECT 31.800 151.100 32.200 153.400 ;
        RECT 33.400 151.100 33.800 153.400 ;
        RECT 36.600 151.100 37.000 153.500 ;
        RECT 39.100 152.800 39.400 153.900 ;
        RECT 41.900 153.800 42.300 153.900 ;
        RECT 45.400 153.600 45.800 155.300 ;
        RECT 47.100 154.200 47.400 155.900 ;
        RECT 47.800 154.800 48.200 155.600 ;
        RECT 48.700 155.200 49.000 155.900 ;
        RECT 51.800 155.800 52.100 157.500 ;
        RECT 53.900 156.400 54.300 157.800 ;
        RECT 53.900 156.100 54.700 156.400 ;
        RECT 51.800 155.500 53.700 155.800 ;
        RECT 50.600 155.200 51.000 155.400 ;
        RECT 48.600 154.900 49.800 155.200 ;
        RECT 50.600 154.900 51.400 155.200 ;
        RECT 48.600 154.800 49.000 154.900 ;
        RECT 47.000 153.800 47.400 154.200 ;
        RECT 43.900 153.300 45.800 153.600 ;
        RECT 43.900 153.200 44.300 153.300 ;
        RECT 45.400 153.100 45.800 153.300 ;
        RECT 46.200 153.100 46.600 153.200 ;
        RECT 47.100 153.100 47.400 153.800 ;
        RECT 48.600 153.100 49.000 153.200 ;
        RECT 49.500 153.100 49.800 154.900 ;
        RECT 51.000 154.800 51.400 154.900 ;
        RECT 50.200 153.800 50.600 154.600 ;
        RECT 51.800 154.400 52.200 155.200 ;
        RECT 52.600 154.400 53.000 155.200 ;
        RECT 53.400 154.500 53.700 155.500 ;
        RECT 53.400 154.100 54.100 154.500 ;
        RECT 54.400 154.200 54.700 156.100 ;
        RECT 55.000 155.100 55.400 155.600 ;
        RECT 56.600 155.100 57.000 159.900 ;
        RECT 55.000 154.800 57.000 155.100 ;
        RECT 53.400 153.900 53.900 154.100 ;
        RECT 45.400 152.800 46.600 153.100 ;
        RECT 47.000 152.800 49.000 153.100 ;
        RECT 38.200 152.100 38.600 152.500 ;
        RECT 39.000 152.400 39.400 152.800 ;
        RECT 39.900 152.700 40.300 152.800 ;
        RECT 39.900 152.400 41.300 152.700 ;
        RECT 41.000 152.100 41.300 152.400 ;
        RECT 43.000 152.100 43.400 152.500 ;
        RECT 38.200 151.800 39.200 152.100 ;
        RECT 38.800 151.100 39.200 151.800 ;
        RECT 41.000 151.100 41.400 152.100 ;
        RECT 43.000 151.800 43.700 152.100 ;
        RECT 43.100 151.100 43.700 151.800 ;
        RECT 45.400 151.100 45.800 152.800 ;
        RECT 46.200 152.400 46.600 152.800 ;
        RECT 47.100 152.100 47.400 152.800 ;
        RECT 48.700 152.400 49.100 152.800 ;
        RECT 47.000 151.100 47.400 152.100 ;
        RECT 49.400 151.100 49.800 153.100 ;
        RECT 51.800 153.600 53.900 153.900 ;
        RECT 54.400 153.800 55.400 154.200 ;
        RECT 51.800 152.500 52.100 153.600 ;
        RECT 54.400 153.500 54.700 153.800 ;
        RECT 54.300 153.300 54.700 153.500 ;
        RECT 53.900 153.000 54.700 153.300 ;
        RECT 51.800 151.500 52.200 152.500 ;
        RECT 53.900 151.500 54.300 153.000 ;
        RECT 56.600 151.100 57.000 154.800 ;
        RECT 57.400 154.100 57.800 154.200 ;
        RECT 58.200 154.100 58.600 154.200 ;
        RECT 57.400 153.800 58.600 154.100 ;
        RECT 57.400 153.200 57.700 153.800 ;
        RECT 58.200 153.400 58.600 153.800 ;
        RECT 57.400 152.400 57.800 153.200 ;
        RECT 59.000 153.100 59.400 159.900 ;
        RECT 60.600 157.500 61.000 159.500 ;
        RECT 59.800 155.800 60.200 156.600 ;
        RECT 60.600 155.800 60.900 157.500 ;
        RECT 62.700 156.400 63.100 159.900 ;
        RECT 62.700 156.100 63.500 156.400 ;
        RECT 60.600 155.500 62.500 155.800 ;
        RECT 60.600 154.400 61.000 155.200 ;
        RECT 61.400 154.400 61.800 155.200 ;
        RECT 62.200 154.500 62.500 155.500 ;
        RECT 62.200 154.100 62.900 154.500 ;
        RECT 63.200 154.200 63.500 156.100 ;
        RECT 63.800 155.100 64.200 155.600 ;
        RECT 65.400 155.100 65.800 159.900 ;
        RECT 63.800 154.800 65.800 155.100 ;
        RECT 63.200 154.100 64.200 154.200 ;
        RECT 64.600 154.100 65.000 154.200 ;
        RECT 62.200 153.900 62.700 154.100 ;
        RECT 60.600 153.600 62.700 153.900 ;
        RECT 63.200 153.800 65.000 154.100 ;
        RECT 59.000 152.800 59.900 153.100 ;
        RECT 59.500 152.200 59.900 152.800 ;
        RECT 59.000 151.800 59.900 152.200 ;
        RECT 59.500 151.100 59.900 151.800 ;
        RECT 60.600 152.500 60.900 153.600 ;
        RECT 63.200 153.500 63.500 153.800 ;
        RECT 63.100 153.300 63.500 153.500 ;
        RECT 62.700 153.000 63.500 153.300 ;
        RECT 60.600 151.500 61.000 152.500 ;
        RECT 62.700 151.500 63.100 153.000 ;
        RECT 65.400 151.100 65.800 154.800 ;
        RECT 67.000 155.600 67.400 159.900 ;
        RECT 69.100 157.900 69.700 159.900 ;
        RECT 71.400 157.900 71.800 159.900 ;
        RECT 73.600 158.200 74.000 159.900 ;
        RECT 73.600 157.900 74.600 158.200 ;
        RECT 69.400 157.500 69.800 157.900 ;
        RECT 71.500 157.600 71.800 157.900 ;
        RECT 71.100 157.300 72.900 157.600 ;
        RECT 74.200 157.500 74.600 157.900 ;
        RECT 71.100 157.200 71.500 157.300 ;
        RECT 72.500 157.200 72.900 157.300 ;
        RECT 69.000 156.600 69.700 157.000 ;
        RECT 69.400 156.100 69.700 156.600 ;
        RECT 70.500 156.500 71.600 156.800 ;
        RECT 70.500 156.400 70.900 156.500 ;
        RECT 69.400 155.800 70.600 156.100 ;
        RECT 67.000 155.300 69.100 155.600 ;
        RECT 67.000 153.600 67.400 155.300 ;
        RECT 68.700 155.200 69.100 155.300 ;
        RECT 70.300 155.200 70.600 155.800 ;
        RECT 71.300 155.900 71.600 156.500 ;
        RECT 71.900 156.500 72.300 156.600 ;
        RECT 74.200 156.500 74.600 156.600 ;
        RECT 71.900 156.200 74.600 156.500 ;
        RECT 71.300 155.700 73.700 155.900 ;
        RECT 75.800 155.700 76.200 159.900 ;
        RECT 76.600 156.200 77.000 159.900 ;
        RECT 78.200 156.200 78.600 159.900 ;
        RECT 76.600 155.900 78.600 156.200 ;
        RECT 79.000 155.900 79.400 159.900 ;
        RECT 71.300 155.600 76.200 155.700 ;
        RECT 73.300 155.500 76.200 155.600 ;
        RECT 73.400 155.400 76.200 155.500 ;
        RECT 77.000 155.200 77.400 155.400 ;
        RECT 79.000 155.200 79.300 155.900 ;
        RECT 79.800 155.700 80.200 159.900 ;
        RECT 82.000 158.200 82.400 159.900 ;
        RECT 81.400 157.900 82.400 158.200 ;
        RECT 84.200 157.900 84.600 159.900 ;
        RECT 86.300 157.900 86.900 159.900 ;
        RECT 81.400 157.500 81.800 157.900 ;
        RECT 84.200 157.600 84.500 157.900 ;
        RECT 83.100 157.300 84.900 157.600 ;
        RECT 86.200 157.500 86.600 157.900 ;
        RECT 83.100 157.200 83.500 157.300 ;
        RECT 84.500 157.200 84.900 157.300 ;
        RECT 81.400 156.500 81.800 156.600 ;
        RECT 83.700 156.500 84.100 156.600 ;
        RECT 81.400 156.200 84.100 156.500 ;
        RECT 84.400 156.500 85.500 156.800 ;
        RECT 84.400 155.900 84.700 156.500 ;
        RECT 85.100 156.400 85.500 156.500 ;
        RECT 86.300 156.600 87.000 157.000 ;
        RECT 86.300 156.100 86.600 156.600 ;
        RECT 82.300 155.700 84.700 155.900 ;
        RECT 79.800 155.600 84.700 155.700 ;
        RECT 85.400 155.800 86.600 156.100 ;
        RECT 79.800 155.500 82.700 155.600 ;
        RECT 79.800 155.400 82.600 155.500 ;
        RECT 67.900 154.900 68.300 155.000 ;
        RECT 67.900 154.600 69.800 154.900 ;
        RECT 70.200 154.800 70.600 155.200 ;
        RECT 72.600 155.100 73.000 155.200 ;
        RECT 72.600 154.800 75.100 155.100 ;
        RECT 76.600 154.900 77.400 155.200 ;
        RECT 78.200 154.900 79.400 155.200 ;
        RECT 83.000 155.100 83.400 155.200 ;
        RECT 76.600 154.800 77.000 154.900 ;
        RECT 69.400 154.500 69.800 154.600 ;
        RECT 70.300 154.200 70.600 154.800 ;
        RECT 74.700 154.700 75.100 154.800 ;
        RECT 73.900 154.200 74.300 154.300 ;
        RECT 70.300 153.900 75.800 154.200 ;
        RECT 70.500 153.800 70.900 153.900 ;
        RECT 67.000 153.300 69.000 153.600 ;
        RECT 66.200 153.100 66.600 153.200 ;
        RECT 67.000 153.100 67.400 153.300 ;
        RECT 68.500 153.200 69.000 153.300 ;
        RECT 66.200 152.800 67.400 153.100 ;
        RECT 68.600 152.800 69.000 153.200 ;
        RECT 73.400 152.800 73.700 153.900 ;
        RECT 75.000 153.800 75.800 153.900 ;
        RECT 77.400 153.800 77.800 154.600 ;
        RECT 66.200 152.400 66.600 152.800 ;
        RECT 67.000 151.100 67.400 152.800 ;
        RECT 72.500 152.700 72.900 152.800 ;
        RECT 69.400 152.100 69.800 152.500 ;
        RECT 71.500 152.400 72.900 152.700 ;
        RECT 73.400 152.400 73.800 152.800 ;
        RECT 71.500 152.100 71.800 152.400 ;
        RECT 74.200 152.100 74.600 152.500 ;
        RECT 69.100 151.800 69.800 152.100 ;
        RECT 69.100 151.100 69.700 151.800 ;
        RECT 71.400 151.100 71.800 152.100 ;
        RECT 73.600 151.800 74.600 152.100 ;
        RECT 73.600 151.100 74.000 151.800 ;
        RECT 75.800 151.100 76.200 153.500 ;
        RECT 78.200 153.100 78.500 154.900 ;
        RECT 79.000 154.800 79.400 154.900 ;
        RECT 80.900 154.800 83.400 155.100 ;
        RECT 79.000 154.200 79.300 154.800 ;
        RECT 80.900 154.700 81.300 154.800 ;
        RECT 82.200 154.700 82.600 154.800 ;
        RECT 81.700 154.200 82.100 154.300 ;
        RECT 85.400 154.200 85.700 155.800 ;
        RECT 88.600 155.600 89.000 159.900 ;
        RECT 86.900 155.300 89.000 155.600 ;
        RECT 91.000 157.500 91.400 159.500 ;
        RECT 93.100 159.200 93.500 159.900 ;
        RECT 92.600 158.800 93.500 159.200 ;
        RECT 91.000 155.800 91.300 157.500 ;
        RECT 93.100 156.400 93.500 158.800 ;
        RECT 93.100 156.100 93.900 156.400 ;
        RECT 91.000 155.500 92.900 155.800 ;
        RECT 86.900 155.200 87.300 155.300 ;
        RECT 87.700 154.900 88.100 155.000 ;
        RECT 86.200 154.600 88.100 154.900 ;
        RECT 86.200 154.500 86.600 154.600 ;
        RECT 79.000 153.800 79.400 154.200 ;
        RECT 80.200 153.900 85.700 154.200 ;
        RECT 80.200 153.800 81.000 153.900 ;
        RECT 78.200 151.100 78.600 153.100 ;
        RECT 79.000 152.800 79.400 153.200 ;
        RECT 78.900 152.400 79.300 152.800 ;
        RECT 79.800 151.100 80.200 153.500 ;
        RECT 82.300 152.800 82.600 153.900 ;
        RECT 85.100 153.800 85.500 153.900 ;
        RECT 88.600 153.600 89.000 155.300 ;
        RECT 91.000 154.400 91.400 155.200 ;
        RECT 91.800 154.400 92.200 155.200 ;
        RECT 92.600 154.500 92.900 155.500 ;
        RECT 92.600 154.100 93.300 154.500 ;
        RECT 93.600 154.200 93.900 156.100 ;
        RECT 94.200 155.100 94.600 155.600 ;
        RECT 95.800 155.100 96.200 159.900 ;
        RECT 94.200 154.800 96.200 155.100 ;
        RECT 92.600 153.900 93.100 154.100 ;
        RECT 87.100 153.300 89.000 153.600 ;
        RECT 87.100 153.200 87.500 153.300 ;
        RECT 81.400 152.100 81.800 152.500 ;
        RECT 82.200 152.400 82.600 152.800 ;
        RECT 83.100 152.700 83.500 152.800 ;
        RECT 83.100 152.400 84.500 152.700 ;
        RECT 84.200 152.100 84.500 152.400 ;
        RECT 86.200 152.100 86.600 152.500 ;
        RECT 81.400 151.800 82.400 152.100 ;
        RECT 82.000 151.100 82.400 151.800 ;
        RECT 84.200 151.100 84.600 152.100 ;
        RECT 86.200 151.800 86.900 152.100 ;
        RECT 86.300 151.100 86.900 151.800 ;
        RECT 88.600 151.100 89.000 153.300 ;
        RECT 91.000 153.600 93.100 153.900 ;
        RECT 93.600 153.800 94.600 154.200 ;
        RECT 91.000 152.500 91.300 153.600 ;
        RECT 93.600 153.500 93.900 153.800 ;
        RECT 93.500 153.300 93.900 153.500 ;
        RECT 93.100 153.000 93.900 153.300 ;
        RECT 91.000 151.500 91.400 152.500 ;
        RECT 93.100 151.500 93.500 153.000 ;
        RECT 95.800 151.100 96.200 154.800 ;
        RECT 98.200 155.100 98.600 159.900 ;
        RECT 100.900 157.200 101.300 159.900 ;
        RECT 103.000 157.500 103.400 159.500 ;
        RECT 100.900 156.800 101.800 157.200 ;
        RECT 100.900 156.400 101.300 156.800 ;
        RECT 100.500 156.100 101.300 156.400 ;
        RECT 99.800 155.100 100.200 155.600 ;
        RECT 98.200 154.800 100.200 155.100 ;
        RECT 96.600 152.400 97.000 153.200 ;
        RECT 97.400 152.400 97.800 153.200 ;
        RECT 98.200 151.100 98.600 154.800 ;
        RECT 100.500 154.200 100.800 156.100 ;
        RECT 103.100 155.800 103.400 157.500 ;
        RECT 101.500 155.500 103.400 155.800 ;
        RECT 103.800 155.600 104.200 159.900 ;
        RECT 105.900 157.900 106.500 159.900 ;
        RECT 108.200 157.900 108.600 159.900 ;
        RECT 110.400 158.200 110.800 159.900 ;
        RECT 110.400 157.900 111.400 158.200 ;
        RECT 106.200 157.500 106.600 157.900 ;
        RECT 108.300 157.600 108.600 157.900 ;
        RECT 107.900 157.300 109.700 157.600 ;
        RECT 111.000 157.500 111.400 157.900 ;
        RECT 107.900 157.200 108.300 157.300 ;
        RECT 109.300 157.200 109.700 157.300 ;
        RECT 105.800 156.600 106.500 157.000 ;
        RECT 106.200 156.100 106.500 156.600 ;
        RECT 107.300 156.500 108.400 156.800 ;
        RECT 107.300 156.400 107.700 156.500 ;
        RECT 106.200 155.800 107.400 156.100 ;
        RECT 101.500 154.500 101.800 155.500 ;
        RECT 103.800 155.300 105.900 155.600 ;
        RECT 99.800 153.800 100.800 154.200 ;
        RECT 101.100 154.100 101.800 154.500 ;
        RECT 102.200 154.400 102.600 155.200 ;
        RECT 103.000 154.400 103.400 155.200 ;
        RECT 100.500 153.500 100.800 153.800 ;
        RECT 101.300 153.900 101.800 154.100 ;
        RECT 101.300 153.600 103.400 153.900 ;
        RECT 100.500 153.300 100.900 153.500 ;
        RECT 100.500 153.000 101.300 153.300 ;
        RECT 100.900 151.500 101.300 153.000 ;
        RECT 103.100 152.500 103.400 153.600 ;
        RECT 103.000 151.500 103.400 152.500 ;
        RECT 103.800 153.600 104.200 155.300 ;
        RECT 105.500 155.200 105.900 155.300 ;
        RECT 104.700 154.900 105.100 155.000 ;
        RECT 104.700 154.600 106.600 154.900 ;
        RECT 106.200 154.500 106.600 154.600 ;
        RECT 107.100 154.200 107.400 155.800 ;
        RECT 108.100 155.900 108.400 156.500 ;
        RECT 108.700 156.500 109.100 156.600 ;
        RECT 111.000 156.500 111.400 156.600 ;
        RECT 108.700 156.200 111.400 156.500 ;
        RECT 108.100 155.700 110.500 155.900 ;
        RECT 112.600 155.700 113.000 159.900 ;
        RECT 108.100 155.600 113.000 155.700 ;
        RECT 110.100 155.500 113.000 155.600 ;
        RECT 110.200 155.400 113.000 155.500 ;
        RECT 113.400 155.600 113.800 159.900 ;
        RECT 115.500 157.900 116.100 159.900 ;
        RECT 117.800 157.900 118.200 159.900 ;
        RECT 120.000 158.200 120.400 159.900 ;
        RECT 120.000 157.900 121.000 158.200 ;
        RECT 115.800 157.500 116.200 157.900 ;
        RECT 117.900 157.600 118.200 157.900 ;
        RECT 117.500 157.300 119.300 157.600 ;
        RECT 120.600 157.500 121.000 157.900 ;
        RECT 117.500 157.200 117.900 157.300 ;
        RECT 118.900 157.200 119.300 157.300 ;
        RECT 115.000 157.000 115.700 157.200 ;
        RECT 115.000 156.800 116.100 157.000 ;
        RECT 115.400 156.600 116.100 156.800 ;
        RECT 115.800 156.100 116.100 156.600 ;
        RECT 116.900 156.500 118.000 156.800 ;
        RECT 116.900 156.400 117.300 156.500 ;
        RECT 115.800 155.800 117.000 156.100 ;
        RECT 113.400 155.300 115.500 155.600 ;
        RECT 109.400 155.100 109.800 155.200 ;
        RECT 109.400 154.800 111.900 155.100 ;
        RECT 111.500 154.700 111.900 154.800 ;
        RECT 110.700 154.200 111.100 154.300 ;
        RECT 107.100 153.900 112.600 154.200 ;
        RECT 107.300 153.800 107.700 153.900 ;
        RECT 103.800 153.300 105.700 153.600 ;
        RECT 103.800 151.100 104.200 153.300 ;
        RECT 105.300 153.200 105.700 153.300 ;
        RECT 110.200 153.200 110.500 153.900 ;
        RECT 111.800 153.800 112.600 153.900 ;
        RECT 113.400 153.600 113.800 155.300 ;
        RECT 115.100 155.200 115.500 155.300 ;
        RECT 114.300 154.900 114.700 155.000 ;
        RECT 114.300 154.600 116.200 154.900 ;
        RECT 115.800 154.500 116.200 154.600 ;
        RECT 116.700 154.200 117.000 155.800 ;
        RECT 117.700 155.900 118.000 156.500 ;
        RECT 118.300 156.500 118.700 156.600 ;
        RECT 120.600 156.500 121.000 156.600 ;
        RECT 118.300 156.200 121.000 156.500 ;
        RECT 117.700 155.700 120.100 155.900 ;
        RECT 122.200 155.700 122.600 159.900 ;
        RECT 117.700 155.600 122.600 155.700 ;
        RECT 119.700 155.500 122.600 155.600 ;
        RECT 119.800 155.400 122.600 155.500 ;
        RECT 119.000 155.100 119.400 155.200 ;
        RECT 123.800 155.100 124.200 159.900 ;
        RECT 126.500 156.400 126.900 159.900 ;
        RECT 128.600 157.500 129.000 159.500 ;
        RECT 126.100 156.100 126.900 156.400 ;
        RECT 125.400 155.100 125.800 155.600 ;
        RECT 119.000 154.800 121.500 155.100 ;
        RECT 121.100 154.700 121.500 154.800 ;
        RECT 123.800 154.800 125.800 155.100 ;
        RECT 120.300 154.200 120.700 154.300 ;
        RECT 116.700 153.900 122.200 154.200 ;
        RECT 116.900 153.800 117.300 153.900 ;
        RECT 119.000 153.800 119.400 153.900 ;
        RECT 109.300 152.700 109.700 152.800 ;
        RECT 106.200 152.100 106.600 152.500 ;
        RECT 108.300 152.400 109.700 152.700 ;
        RECT 110.200 152.400 110.600 153.200 ;
        RECT 108.300 152.100 108.600 152.400 ;
        RECT 111.000 152.100 111.400 152.500 ;
        RECT 105.900 151.800 106.600 152.100 ;
        RECT 105.900 151.100 106.500 151.800 ;
        RECT 108.200 151.100 108.600 152.100 ;
        RECT 110.400 151.800 111.400 152.100 ;
        RECT 110.400 151.100 110.800 151.800 ;
        RECT 112.600 151.100 113.000 153.500 ;
        RECT 113.400 153.300 115.300 153.600 ;
        RECT 113.400 151.100 113.800 153.300 ;
        RECT 114.900 153.200 115.300 153.300 ;
        RECT 119.800 152.800 120.100 153.900 ;
        RECT 121.400 153.800 122.200 153.900 ;
        RECT 118.900 152.700 119.300 152.800 ;
        RECT 115.800 152.100 116.200 152.500 ;
        RECT 117.900 152.400 119.300 152.700 ;
        RECT 119.800 152.400 120.200 152.800 ;
        RECT 117.900 152.100 118.200 152.400 ;
        RECT 120.600 152.100 121.000 152.500 ;
        RECT 115.500 151.800 116.200 152.100 ;
        RECT 115.500 151.100 116.100 151.800 ;
        RECT 117.800 151.100 118.200 152.100 ;
        RECT 120.000 151.800 121.000 152.100 ;
        RECT 120.000 151.100 120.400 151.800 ;
        RECT 122.200 151.100 122.600 153.500 ;
        RECT 123.000 152.400 123.400 153.200 ;
        RECT 123.800 151.100 124.200 154.800 ;
        RECT 126.100 154.200 126.400 156.100 ;
        RECT 128.700 155.800 129.000 157.500 ;
        RECT 127.100 155.500 129.000 155.800 ;
        RECT 129.400 157.500 129.800 159.500 ;
        RECT 129.400 155.800 129.700 157.500 ;
        RECT 131.500 156.400 131.900 159.900 ;
        RECT 131.500 156.100 132.300 156.400 ;
        RECT 129.400 155.500 131.300 155.800 ;
        RECT 127.100 154.500 127.400 155.500 ;
        RECT 125.400 153.800 126.400 154.200 ;
        RECT 126.700 154.100 127.400 154.500 ;
        RECT 127.800 154.400 128.200 155.200 ;
        RECT 128.600 154.400 129.000 155.200 ;
        RECT 129.400 154.400 129.800 155.200 ;
        RECT 130.200 154.400 130.600 155.200 ;
        RECT 131.000 154.500 131.300 155.500 ;
        RECT 126.100 153.500 126.400 153.800 ;
        RECT 126.900 153.900 127.400 154.100 ;
        RECT 131.000 154.100 131.700 154.500 ;
        RECT 132.000 154.200 132.300 156.100 ;
        RECT 132.600 155.100 133.000 155.600 ;
        RECT 134.200 155.100 134.600 159.900 ;
        RECT 137.400 155.700 137.800 159.900 ;
        RECT 139.600 158.200 140.000 159.900 ;
        RECT 139.000 157.900 140.000 158.200 ;
        RECT 141.800 157.900 142.200 159.900 ;
        RECT 143.900 157.900 144.500 159.900 ;
        RECT 139.000 157.500 139.400 157.900 ;
        RECT 141.800 157.600 142.100 157.900 ;
        RECT 140.700 157.300 142.500 157.600 ;
        RECT 143.800 157.500 144.200 157.900 ;
        RECT 140.700 157.200 141.100 157.300 ;
        RECT 142.100 157.200 142.500 157.300 ;
        RECT 139.000 156.500 139.400 156.600 ;
        RECT 141.300 156.500 141.700 156.600 ;
        RECT 139.000 156.200 141.700 156.500 ;
        RECT 142.000 156.500 143.100 156.800 ;
        RECT 142.000 155.900 142.300 156.500 ;
        RECT 142.700 156.400 143.100 156.500 ;
        RECT 143.900 156.600 144.600 157.000 ;
        RECT 143.900 156.100 144.200 156.600 ;
        RECT 139.900 155.700 142.300 155.900 ;
        RECT 137.400 155.600 142.300 155.700 ;
        RECT 143.000 155.800 144.200 156.100 ;
        RECT 137.400 155.500 140.300 155.600 ;
        RECT 137.400 155.400 140.200 155.500 ;
        RECT 140.600 155.100 141.000 155.200 ;
        RECT 132.600 154.800 134.600 155.100 ;
        RECT 132.000 154.100 133.000 154.200 ;
        RECT 133.400 154.100 133.800 154.200 ;
        RECT 131.000 153.900 131.500 154.100 ;
        RECT 126.900 153.600 129.000 153.900 ;
        RECT 126.100 153.300 126.500 153.500 ;
        RECT 126.100 153.000 126.900 153.300 ;
        RECT 126.500 151.500 126.900 153.000 ;
        RECT 128.700 152.500 129.000 153.600 ;
        RECT 128.600 151.500 129.000 152.500 ;
        RECT 129.400 153.600 131.500 153.900 ;
        RECT 132.000 153.800 133.800 154.100 ;
        RECT 129.400 152.500 129.700 153.600 ;
        RECT 132.000 153.500 132.300 153.800 ;
        RECT 131.900 153.300 132.300 153.500 ;
        RECT 131.500 153.000 132.300 153.300 ;
        RECT 129.400 151.500 129.800 152.500 ;
        RECT 131.500 151.500 131.900 153.000 ;
        RECT 134.200 151.100 134.600 154.800 ;
        RECT 138.500 154.800 141.000 155.100 ;
        RECT 138.500 154.700 138.900 154.800 ;
        RECT 139.800 154.700 140.200 154.800 ;
        RECT 139.300 154.200 139.700 154.300 ;
        RECT 143.000 154.200 143.300 155.800 ;
        RECT 146.200 155.600 146.600 159.900 ;
        RECT 144.500 155.300 146.600 155.600 ;
        RECT 144.500 155.200 144.900 155.300 ;
        RECT 145.300 154.900 145.700 155.000 ;
        RECT 143.800 154.600 145.700 154.900 ;
        RECT 143.800 154.500 144.200 154.600 ;
        RECT 137.800 153.900 143.300 154.200 ;
        RECT 137.800 153.800 138.600 153.900 ;
        RECT 135.000 152.400 135.400 153.200 ;
        RECT 137.400 151.100 137.800 153.500 ;
        RECT 139.900 153.200 140.200 153.900 ;
        RECT 142.700 153.800 143.100 153.900 ;
        RECT 146.200 153.600 146.600 155.300 ;
        RECT 147.800 155.600 148.200 159.900 ;
        RECT 149.400 155.600 149.800 159.900 ;
        RECT 151.000 155.600 151.400 159.900 ;
        RECT 152.600 155.600 153.000 159.900 ;
        RECT 147.800 155.200 148.700 155.600 ;
        RECT 149.400 155.200 150.500 155.600 ;
        RECT 151.000 155.200 152.100 155.600 ;
        RECT 152.600 155.200 153.800 155.600 ;
        RECT 148.300 154.500 148.700 155.200 ;
        RECT 150.100 154.500 150.500 155.200 ;
        RECT 151.700 154.500 152.100 155.200 ;
        RECT 148.300 154.100 149.600 154.500 ;
        RECT 150.100 154.100 151.300 154.500 ;
        RECT 151.700 154.100 153.000 154.500 ;
        RECT 148.300 153.800 148.700 154.100 ;
        RECT 150.100 153.800 150.500 154.100 ;
        RECT 151.700 153.800 152.100 154.100 ;
        RECT 153.400 153.800 153.800 155.200 ;
        RECT 144.700 153.300 146.600 153.600 ;
        RECT 144.700 153.200 145.100 153.300 ;
        RECT 139.000 152.100 139.400 152.500 ;
        RECT 139.800 152.400 140.200 153.200 ;
        RECT 140.700 152.700 141.100 152.800 ;
        RECT 140.700 152.400 142.100 152.700 ;
        RECT 141.800 152.100 142.100 152.400 ;
        RECT 143.800 152.100 144.200 152.500 ;
        RECT 139.000 151.800 140.000 152.100 ;
        RECT 139.600 151.100 140.000 151.800 ;
        RECT 141.800 151.100 142.200 152.100 ;
        RECT 143.800 151.800 144.500 152.100 ;
        RECT 143.900 151.100 144.500 151.800 ;
        RECT 146.200 151.100 146.600 153.300 ;
        RECT 147.800 153.400 148.700 153.800 ;
        RECT 149.400 153.400 150.500 153.800 ;
        RECT 151.000 153.400 152.100 153.800 ;
        RECT 152.600 153.400 153.800 153.800 ;
        RECT 147.800 151.100 148.200 153.400 ;
        RECT 149.400 151.100 149.800 153.400 ;
        RECT 151.000 151.100 151.400 153.400 ;
        RECT 152.600 151.100 153.000 153.400 ;
        RECT 154.200 152.400 154.600 153.200 ;
        RECT 155.000 151.100 155.400 159.900 ;
        RECT 156.600 158.200 157.000 159.900 ;
        RECT 156.500 157.900 157.000 158.200 ;
        RECT 156.500 157.600 156.800 157.900 ;
        RECT 158.200 157.600 158.600 159.900 ;
        RECT 159.800 158.500 160.200 159.900 ;
        RECT 160.600 158.500 161.000 159.900 ;
        RECT 155.800 157.300 156.800 157.600 ;
        RECT 155.800 154.500 156.200 157.300 ;
        RECT 157.100 157.200 159.200 157.600 ;
        RECT 161.400 157.500 161.800 159.900 ;
        RECT 163.000 157.500 163.400 159.900 ;
        RECT 157.100 157.000 157.400 157.200 ;
        RECT 156.600 156.600 157.400 157.000 ;
        RECT 158.900 156.900 161.800 157.200 ;
        RECT 157.900 156.600 158.600 156.900 ;
        RECT 157.900 156.500 161.000 156.600 ;
        RECT 158.300 156.300 161.000 156.500 ;
        RECT 160.600 156.200 161.000 156.300 ;
        RECT 161.500 156.500 161.800 156.900 ;
        RECT 162.100 156.800 163.400 157.200 ;
        RECT 164.600 156.800 165.000 159.900 ;
        RECT 165.400 158.500 165.800 159.900 ;
        RECT 166.200 158.500 166.600 159.900 ;
        RECT 167.000 158.500 167.400 159.900 ;
        RECT 166.200 157.200 168.300 157.600 ;
        RECT 168.600 157.200 169.000 159.900 ;
        RECT 170.200 157.600 170.600 159.900 ;
        RECT 170.200 157.300 171.500 157.600 ;
        RECT 168.600 156.800 169.900 157.200 ;
        RECT 165.400 156.500 165.800 156.600 ;
        RECT 161.500 156.200 165.800 156.500 ;
        RECT 167.000 156.500 167.400 156.600 ;
        RECT 171.200 156.500 171.500 157.300 ;
        RECT 167.000 156.200 171.500 156.500 ;
        RECT 171.200 155.300 171.500 156.200 ;
        RECT 171.800 156.000 172.200 159.900 ;
        RECT 173.400 156.200 173.800 159.900 ;
        RECT 171.800 155.600 172.300 156.000 ;
        RECT 173.400 155.900 174.500 156.200 ;
        RECT 171.200 155.000 171.600 155.300 ;
        RECT 155.800 154.100 160.200 154.500 ;
        RECT 160.500 154.300 161.500 154.700 ;
        RECT 163.400 154.300 165.000 154.700 ;
        RECT 155.800 151.100 156.200 154.100 ;
        RECT 157.000 153.400 158.500 153.800 ;
        RECT 158.100 153.100 158.500 153.400 ;
        RECT 161.100 153.100 161.500 154.300 ;
        RECT 162.200 153.400 162.600 154.200 ;
        RECT 164.800 153.900 165.200 154.000 ;
        RECT 163.000 153.600 165.200 153.900 ;
        RECT 163.000 153.500 163.400 153.600 ;
        RECT 166.200 153.200 166.600 154.600 ;
        RECT 169.100 154.300 171.000 154.700 ;
        RECT 169.100 153.700 169.500 154.300 ;
        RECT 171.300 154.000 171.600 155.000 ;
        RECT 163.000 153.100 163.400 153.200 ;
        RECT 158.100 152.700 159.400 153.100 ;
        RECT 161.100 152.800 163.400 153.100 ;
        RECT 163.800 152.800 164.600 153.200 ;
        RECT 166.100 152.800 166.600 153.200 ;
        RECT 168.600 153.400 169.500 153.700 ;
        RECT 171.000 153.700 171.600 154.000 ;
        RECT 168.600 153.100 169.000 153.400 ;
        RECT 159.000 151.100 159.400 152.700 ;
        RECT 167.800 152.700 169.000 153.100 ;
        RECT 159.800 151.100 160.200 152.500 ;
        RECT 160.600 151.100 161.000 152.500 ;
        RECT 161.400 151.100 161.800 152.500 ;
        RECT 163.000 151.100 163.400 152.500 ;
        RECT 164.600 151.100 165.000 152.500 ;
        RECT 165.400 151.100 165.800 152.500 ;
        RECT 166.200 151.100 166.600 152.500 ;
        RECT 167.000 151.100 167.400 152.500 ;
        RECT 167.800 151.100 168.200 152.700 ;
        RECT 171.000 151.100 171.400 153.700 ;
        RECT 171.900 153.400 172.300 155.600 ;
        RECT 174.200 155.600 174.500 155.900 ;
        RECT 174.200 155.200 174.800 155.600 ;
        RECT 173.400 154.400 173.800 155.200 ;
        RECT 174.200 153.700 174.500 155.200 ;
        RECT 171.800 153.000 172.300 153.400 ;
        RECT 173.400 153.400 174.500 153.700 ;
        RECT 171.800 151.100 172.200 153.000 ;
        RECT 173.400 151.100 173.800 153.400 ;
        RECT 175.800 151.100 176.200 159.900 ;
        RECT 177.400 156.200 177.800 159.900 ;
        RECT 177.400 155.900 178.500 156.200 ;
        RECT 178.200 155.600 178.500 155.900 ;
        RECT 178.200 155.200 178.800 155.600 ;
        RECT 177.400 154.400 177.800 155.200 ;
        RECT 178.200 153.700 178.500 155.200 ;
        RECT 177.400 153.400 178.500 153.700 ;
        RECT 176.600 152.400 177.000 153.200 ;
        RECT 177.400 151.100 177.800 153.400 ;
        RECT 0.600 147.500 1.000 149.900 ;
        RECT 2.800 149.200 3.200 149.900 ;
        RECT 2.200 148.900 3.200 149.200 ;
        RECT 5.000 148.900 5.400 149.900 ;
        RECT 7.100 149.200 7.700 149.900 ;
        RECT 7.000 148.900 7.700 149.200 ;
        RECT 2.200 148.500 2.600 148.900 ;
        RECT 5.000 148.600 5.300 148.900 ;
        RECT 3.000 148.200 3.400 148.600 ;
        RECT 3.900 148.300 5.300 148.600 ;
        RECT 7.000 148.500 7.400 148.900 ;
        RECT 3.900 148.200 4.300 148.300 ;
        RECT 1.000 147.100 1.800 147.200 ;
        RECT 3.100 147.100 3.400 148.200 ;
        RECT 7.900 147.700 8.300 147.800 ;
        RECT 9.400 147.700 9.800 149.900 ;
        RECT 11.000 148.900 11.400 149.900 ;
        RECT 10.200 147.800 10.600 148.600 ;
        RECT 11.100 148.100 11.400 148.900 ;
        RECT 12.700 148.200 13.100 148.600 ;
        RECT 12.600 148.100 13.000 148.200 ;
        RECT 11.000 147.800 13.000 148.100 ;
        RECT 13.400 147.900 13.800 149.900 ;
        RECT 17.100 148.200 17.500 149.900 ;
        RECT 7.900 147.400 9.800 147.700 ;
        RECT 5.900 147.100 6.300 147.200 ;
        RECT 1.000 146.800 6.500 147.100 ;
        RECT 2.500 146.700 2.900 146.800 ;
        RECT 1.700 146.200 2.100 146.300 ;
        RECT 6.200 146.200 6.500 146.800 ;
        RECT 7.000 146.400 7.400 146.500 ;
        RECT 1.700 145.900 4.200 146.200 ;
        RECT 3.800 145.800 4.200 145.900 ;
        RECT 6.200 145.800 6.600 146.200 ;
        RECT 7.000 146.100 8.900 146.400 ;
        RECT 8.500 146.000 8.900 146.100 ;
        RECT 0.600 145.500 3.400 145.600 ;
        RECT 0.600 145.400 3.500 145.500 ;
        RECT 0.600 145.300 5.500 145.400 ;
        RECT 0.600 141.100 1.000 145.300 ;
        RECT 3.100 145.100 5.500 145.300 ;
        RECT 2.200 144.500 4.900 144.800 ;
        RECT 2.200 144.400 2.600 144.500 ;
        RECT 4.500 144.400 4.900 144.500 ;
        RECT 5.200 144.500 5.500 145.100 ;
        RECT 6.200 145.200 6.500 145.800 ;
        RECT 7.700 145.700 8.100 145.800 ;
        RECT 9.400 145.700 9.800 147.400 ;
        RECT 11.100 147.200 11.400 147.800 ;
        RECT 11.000 146.800 11.400 147.200 ;
        RECT 7.700 145.400 9.800 145.700 ;
        RECT 6.200 144.900 7.400 145.200 ;
        RECT 5.900 144.500 6.300 144.600 ;
        RECT 5.200 144.200 6.300 144.500 ;
        RECT 7.100 144.400 7.400 144.900 ;
        RECT 7.100 144.000 7.800 144.400 ;
        RECT 3.900 143.700 4.300 143.800 ;
        RECT 5.300 143.700 5.700 143.800 ;
        RECT 2.200 143.100 2.600 143.500 ;
        RECT 3.900 143.400 5.700 143.700 ;
        RECT 5.000 143.100 5.300 143.400 ;
        RECT 7.000 143.100 7.400 143.500 ;
        RECT 2.200 142.800 3.200 143.100 ;
        RECT 2.800 141.100 3.200 142.800 ;
        RECT 5.000 141.100 5.400 143.100 ;
        RECT 7.100 141.100 7.700 143.100 ;
        RECT 9.400 141.100 9.800 145.400 ;
        RECT 11.100 145.100 11.400 146.800 ;
        RECT 12.600 146.800 13.000 147.200 ;
        RECT 12.600 146.200 12.900 146.800 ;
        RECT 11.800 145.400 12.200 146.200 ;
        RECT 12.600 146.100 13.000 146.200 ;
        RECT 13.500 146.100 13.800 147.900 ;
        RECT 16.600 147.900 17.500 148.200 ;
        RECT 20.000 148.200 20.400 149.900 ;
        RECT 21.400 148.500 21.800 149.500 ;
        RECT 14.200 146.400 14.600 147.200 ;
        RECT 15.800 146.800 16.200 147.600 ;
        RECT 15.000 146.100 15.400 146.200 ;
        RECT 12.600 145.800 13.800 146.100 ;
        RECT 14.600 145.800 15.400 146.100 ;
        RECT 16.600 146.100 17.000 147.900 ;
        RECT 20.000 147.800 21.000 148.200 ;
        RECT 20.000 147.100 20.400 147.800 ;
        RECT 21.400 147.400 21.700 148.500 ;
        RECT 23.500 148.000 23.900 149.500 ;
        RECT 23.500 147.700 24.300 148.000 ;
        RECT 23.900 147.500 24.300 147.700 ;
        RECT 21.400 147.100 23.500 147.400 ;
        RECT 20.000 146.900 20.900 147.100 ;
        RECT 20.100 146.800 20.900 146.900 ;
        RECT 16.600 145.800 18.600 146.100 ;
        RECT 19.000 145.800 19.800 146.200 ;
        RECT 12.700 145.100 13.000 145.800 ;
        RECT 14.600 145.600 15.000 145.800 ;
        RECT 11.000 144.700 11.900 145.100 ;
        RECT 11.500 141.100 11.900 144.700 ;
        RECT 12.600 141.100 13.000 145.100 ;
        RECT 13.400 144.800 15.400 145.100 ;
        RECT 13.400 141.100 13.800 144.800 ;
        RECT 15.000 141.100 15.400 144.800 ;
        RECT 16.600 141.100 17.000 145.800 ;
        RECT 17.400 144.400 17.800 145.200 ;
        RECT 18.200 144.800 18.600 145.800 ;
        RECT 20.600 145.200 20.900 146.800 ;
        RECT 23.000 146.900 23.500 147.100 ;
        RECT 24.000 147.200 24.300 147.500 ;
        RECT 24.000 147.100 25.000 147.200 ;
        RECT 25.400 147.100 25.800 147.200 ;
        RECT 21.400 145.800 21.800 146.600 ;
        RECT 22.200 145.800 22.600 146.600 ;
        RECT 23.000 146.500 23.700 146.900 ;
        RECT 24.000 146.800 25.800 147.100 ;
        RECT 23.000 145.500 23.300 146.500 ;
        RECT 21.400 145.200 23.300 145.500 ;
        RECT 20.600 144.800 21.000 145.200 ;
        RECT 18.200 144.100 18.600 144.200 ;
        RECT 19.800 144.100 20.200 144.600 ;
        RECT 18.200 143.800 20.200 144.100 ;
        RECT 20.600 143.500 20.900 144.800 ;
        RECT 19.100 143.200 20.900 143.500 ;
        RECT 19.100 143.100 19.400 143.200 ;
        RECT 19.000 141.100 19.400 143.100 ;
        RECT 20.600 143.100 20.900 143.200 ;
        RECT 21.400 143.500 21.700 145.200 ;
        RECT 24.000 144.900 24.300 146.800 ;
        RECT 24.600 146.100 25.000 146.200 ;
        RECT 26.200 146.100 26.600 149.900 ;
        RECT 27.000 148.100 27.400 148.600 ;
        RECT 27.800 148.100 28.200 149.900 ;
        RECT 29.900 149.200 30.500 149.900 ;
        RECT 29.900 148.900 30.600 149.200 ;
        RECT 32.200 148.900 32.600 149.900 ;
        RECT 34.400 149.200 34.800 149.900 ;
        RECT 34.400 148.900 35.400 149.200 ;
        RECT 30.200 148.500 30.600 148.900 ;
        RECT 32.300 148.600 32.600 148.900 ;
        RECT 32.300 148.300 33.700 148.600 ;
        RECT 33.300 148.200 33.700 148.300 ;
        RECT 34.200 148.200 34.600 148.600 ;
        RECT 35.000 148.500 35.400 148.900 ;
        RECT 27.000 147.800 28.200 148.100 ;
        RECT 24.600 145.800 26.600 146.100 ;
        RECT 24.600 145.400 25.000 145.800 ;
        RECT 23.500 144.600 24.300 144.900 ;
        RECT 20.600 141.100 21.000 143.100 ;
        RECT 21.400 141.500 21.800 143.500 ;
        RECT 23.500 141.100 23.900 144.600 ;
        RECT 26.200 141.100 26.600 145.800 ;
        RECT 27.800 147.700 28.200 147.800 ;
        RECT 29.300 147.700 29.700 147.800 ;
        RECT 27.800 147.400 29.700 147.700 ;
        RECT 27.800 145.700 28.200 147.400 ;
        RECT 31.300 147.100 31.700 147.200 ;
        RECT 34.200 147.100 34.500 148.200 ;
        RECT 36.600 147.500 37.000 149.900 ;
        RECT 40.600 147.900 41.000 149.900 ;
        RECT 43.000 148.900 43.400 149.900 ;
        RECT 41.300 148.200 41.700 148.600 ;
        RECT 41.400 148.100 41.800 148.200 ;
        RECT 43.000 148.100 43.300 148.900 ;
        RECT 35.800 147.100 36.600 147.200 ;
        RECT 31.100 146.800 36.600 147.100 ;
        RECT 30.200 146.400 30.600 146.500 ;
        RECT 28.700 146.100 30.600 146.400 ;
        RECT 28.700 146.000 29.100 146.100 ;
        RECT 29.500 145.700 29.900 145.800 ;
        RECT 27.800 145.400 29.900 145.700 ;
        RECT 27.800 141.100 28.200 145.400 ;
        RECT 31.100 145.200 31.400 146.800 ;
        RECT 34.700 146.700 35.100 146.800 ;
        RECT 39.800 146.400 40.200 147.200 ;
        RECT 35.500 146.200 35.900 146.300 ;
        RECT 33.400 145.900 35.900 146.200 ;
        RECT 39.000 146.100 39.400 146.200 ;
        RECT 40.600 146.100 40.900 147.900 ;
        RECT 41.400 147.800 43.300 148.100 ;
        RECT 43.800 147.800 44.200 148.600 ;
        RECT 45.900 148.200 46.300 149.900 ;
        RECT 45.400 147.900 46.300 148.200 ;
        RECT 43.000 147.200 43.300 147.800 ;
        RECT 43.000 146.800 43.400 147.200 ;
        RECT 44.600 146.800 45.000 147.600 ;
        RECT 41.400 146.100 41.800 146.200 ;
        RECT 33.400 145.800 33.800 145.900 ;
        RECT 39.000 145.800 39.800 146.100 ;
        RECT 40.600 145.800 41.800 146.100 ;
        RECT 39.400 145.600 39.800 145.800 ;
        RECT 34.200 145.500 37.000 145.600 ;
        RECT 34.100 145.400 37.000 145.500 ;
        RECT 30.200 144.900 31.400 145.200 ;
        RECT 32.100 145.300 37.000 145.400 ;
        RECT 32.100 145.100 34.500 145.300 ;
        RECT 30.200 144.400 30.500 144.900 ;
        RECT 29.800 144.000 30.500 144.400 ;
        RECT 31.300 144.500 31.700 144.600 ;
        RECT 32.100 144.500 32.400 145.100 ;
        RECT 31.300 144.200 32.400 144.500 ;
        RECT 32.700 144.500 35.400 144.800 ;
        RECT 32.700 144.400 33.100 144.500 ;
        RECT 35.000 144.400 35.400 144.500 ;
        RECT 31.900 143.700 32.300 143.800 ;
        RECT 33.300 143.700 33.700 143.800 ;
        RECT 30.200 143.100 30.600 143.500 ;
        RECT 31.900 143.400 33.700 143.700 ;
        RECT 32.300 143.100 32.600 143.400 ;
        RECT 35.000 143.100 35.400 143.500 ;
        RECT 29.900 141.100 30.500 143.100 ;
        RECT 32.200 141.100 32.600 143.100 ;
        RECT 34.400 142.800 35.400 143.100 ;
        RECT 34.400 141.100 34.800 142.800 ;
        RECT 36.600 141.100 37.000 145.300 ;
        RECT 41.400 145.200 41.700 145.800 ;
        RECT 42.200 145.400 42.600 146.200 ;
        RECT 39.000 144.800 41.000 145.100 ;
        RECT 39.000 141.100 39.400 144.800 ;
        RECT 40.600 141.100 41.000 144.800 ;
        RECT 41.400 141.100 41.800 145.200 ;
        RECT 43.000 145.100 43.300 146.800 ;
        RECT 42.500 144.700 43.400 145.100 ;
        RECT 42.500 141.100 42.900 144.700 ;
        RECT 45.400 141.100 45.800 147.900 ;
        RECT 47.000 147.500 47.400 149.900 ;
        RECT 49.200 149.200 49.600 149.900 ;
        RECT 48.600 148.900 49.600 149.200 ;
        RECT 51.400 148.900 51.800 149.900 ;
        RECT 53.500 149.200 54.100 149.900 ;
        RECT 53.400 148.900 54.100 149.200 ;
        RECT 48.600 148.500 49.000 148.900 ;
        RECT 51.400 148.600 51.700 148.900 ;
        RECT 49.400 147.800 49.800 148.600 ;
        RECT 50.300 148.300 51.700 148.600 ;
        RECT 53.400 148.500 53.800 148.900 ;
        RECT 50.300 148.200 50.700 148.300 ;
        RECT 47.400 147.100 48.200 147.200 ;
        RECT 49.500 147.100 49.800 147.800 ;
        RECT 54.300 147.700 54.700 147.800 ;
        RECT 55.800 147.700 56.200 149.900 ;
        RECT 54.300 147.400 56.200 147.700 ;
        RECT 52.300 147.100 52.700 147.200 ;
        RECT 47.400 146.800 52.900 147.100 ;
        RECT 48.900 146.700 49.300 146.800 ;
        RECT 48.100 146.200 48.500 146.300 ;
        RECT 49.400 146.200 49.800 146.300 ;
        RECT 48.100 145.900 50.600 146.200 ;
        RECT 50.200 145.800 50.600 145.900 ;
        RECT 47.000 145.500 49.800 145.600 ;
        RECT 47.000 145.400 49.900 145.500 ;
        RECT 47.000 145.300 51.900 145.400 ;
        RECT 46.200 144.400 46.600 145.200 ;
        RECT 47.000 141.100 47.400 145.300 ;
        RECT 49.500 145.100 51.900 145.300 ;
        RECT 48.600 144.500 51.300 144.800 ;
        RECT 48.600 144.400 49.000 144.500 ;
        RECT 50.900 144.400 51.300 144.500 ;
        RECT 51.600 144.500 51.900 145.100 ;
        RECT 52.600 145.200 52.900 146.800 ;
        RECT 53.400 146.400 53.800 146.500 ;
        RECT 53.400 146.100 55.300 146.400 ;
        RECT 54.900 146.000 55.300 146.100 ;
        RECT 54.100 145.700 54.500 145.800 ;
        RECT 55.800 145.700 56.200 147.400 ;
        RECT 57.200 147.100 57.600 149.900 ;
        RECT 61.100 148.200 61.500 149.900 ;
        RECT 63.800 149.200 64.200 149.900 ;
        RECT 63.800 148.900 64.300 149.200 ;
        RECT 64.000 148.800 64.300 148.900 ;
        RECT 65.400 148.900 65.800 149.900 ;
        RECT 67.800 149.100 68.200 149.200 ;
        RECT 68.600 149.100 69.000 149.900 ;
        RECT 65.400 148.800 66.000 148.900 ;
        RECT 67.800 148.800 69.000 149.100 ;
        RECT 70.700 149.200 71.300 149.900 ;
        RECT 70.700 148.900 71.400 149.200 ;
        RECT 73.000 148.900 73.400 149.900 ;
        RECT 75.200 149.200 75.600 149.900 ;
        RECT 75.200 148.900 76.200 149.200 ;
        RECT 64.000 148.500 66.000 148.800 ;
        RECT 60.600 147.900 61.500 148.200 ;
        RECT 54.100 145.400 56.200 145.700 ;
        RECT 52.600 144.900 53.800 145.200 ;
        RECT 52.300 144.500 52.700 144.600 ;
        RECT 51.600 144.200 52.700 144.500 ;
        RECT 53.500 144.400 53.800 144.900 ;
        RECT 53.500 144.000 54.200 144.400 ;
        RECT 50.300 143.700 50.700 143.800 ;
        RECT 51.700 143.700 52.100 143.800 ;
        RECT 48.600 143.100 49.000 143.500 ;
        RECT 50.300 143.400 52.100 143.700 ;
        RECT 51.400 143.100 51.700 143.400 ;
        RECT 53.400 143.100 53.800 143.500 ;
        RECT 48.600 142.800 49.600 143.100 ;
        RECT 49.200 141.100 49.600 142.800 ;
        RECT 51.400 141.100 51.800 143.100 ;
        RECT 53.500 141.100 54.100 143.100 ;
        RECT 55.800 141.100 56.200 145.400 ;
        RECT 56.700 146.900 57.600 147.100 ;
        RECT 56.700 146.800 57.500 146.900 ;
        RECT 59.800 146.800 60.200 147.600 ;
        RECT 56.700 145.200 57.000 146.800 ;
        RECT 57.400 145.800 58.600 146.200 ;
        RECT 56.600 144.800 57.000 145.200 ;
        RECT 59.000 145.100 59.400 145.600 ;
        RECT 60.600 145.100 61.000 147.900 ;
        RECT 63.000 147.800 63.900 148.200 ;
        RECT 63.800 146.800 64.600 147.200 ;
        RECT 65.700 147.100 66.000 148.500 ;
        RECT 68.600 147.700 69.000 148.800 ;
        RECT 71.000 148.500 71.400 148.900 ;
        RECT 73.100 148.600 73.400 148.900 ;
        RECT 73.100 148.300 74.500 148.600 ;
        RECT 74.100 148.200 74.500 148.300 ;
        RECT 75.000 147.800 75.400 148.600 ;
        RECT 75.800 148.500 76.200 148.900 ;
        RECT 70.100 147.700 70.500 147.800 ;
        RECT 68.600 147.400 70.500 147.700 ;
        RECT 67.000 147.100 67.400 147.200 ;
        RECT 65.700 146.800 67.400 147.100 ;
        RECT 64.600 145.800 65.400 146.200 ;
        RECT 65.700 145.200 66.000 146.800 ;
        RECT 68.600 145.700 69.000 147.400 ;
        RECT 72.100 147.100 72.500 147.200 ;
        RECT 75.000 147.100 75.300 147.800 ;
        RECT 77.400 147.500 77.800 149.900 ;
        RECT 79.000 148.800 79.400 149.900 ;
        RECT 79.000 147.200 79.300 148.800 ;
        RECT 79.800 147.800 80.200 148.600 ;
        RECT 80.600 148.500 81.000 149.500 ;
        RECT 80.600 147.400 80.900 148.500 ;
        RECT 82.700 148.000 83.100 149.500 ;
        RECT 82.700 147.700 83.500 148.000 ;
        RECT 83.100 147.500 83.500 147.700 ;
        RECT 76.600 147.100 77.400 147.200 ;
        RECT 71.900 146.800 77.400 147.100 ;
        RECT 79.000 146.800 79.400 147.200 ;
        RECT 80.600 147.100 82.700 147.400 ;
        RECT 82.200 146.900 82.700 147.100 ;
        RECT 83.200 147.200 83.500 147.500 ;
        RECT 83.200 147.100 84.200 147.200 ;
        RECT 84.600 147.100 85.000 147.200 ;
        RECT 71.000 146.400 71.400 146.500 ;
        RECT 69.500 146.100 71.400 146.400 ;
        RECT 69.500 146.000 69.900 146.100 ;
        RECT 70.300 145.700 70.700 145.800 ;
        RECT 68.600 145.400 70.700 145.700 ;
        RECT 59.000 144.800 61.000 145.100 ;
        RECT 56.700 143.500 57.000 144.800 ;
        RECT 57.400 144.100 57.800 144.600 ;
        RECT 59.000 144.100 59.400 144.200 ;
        RECT 57.400 143.800 59.400 144.100 ;
        RECT 56.700 143.200 58.500 143.500 ;
        RECT 56.700 143.100 57.000 143.200 ;
        RECT 56.600 141.100 57.000 143.100 ;
        RECT 58.200 143.100 58.500 143.200 ;
        RECT 58.200 141.100 58.600 143.100 ;
        RECT 60.600 141.100 61.000 144.800 ;
        RECT 61.400 144.400 61.800 145.200 ;
        RECT 65.700 144.900 67.400 145.200 ;
        RECT 67.000 144.800 67.400 144.900 ;
        RECT 62.300 144.400 64.100 144.700 ;
        RECT 62.300 144.100 62.600 144.400 ;
        RECT 62.200 141.100 62.600 144.100 ;
        RECT 63.800 144.100 64.100 144.400 ;
        RECT 64.700 144.500 66.500 144.600 ;
        RECT 67.000 144.500 67.300 144.800 ;
        RECT 64.700 144.300 66.600 144.500 ;
        RECT 64.700 144.100 65.000 144.300 ;
        RECT 63.800 141.400 64.200 144.100 ;
        RECT 64.600 141.700 65.000 144.100 ;
        RECT 65.400 141.400 65.800 144.000 ;
        RECT 66.200 141.500 66.600 144.300 ;
        RECT 67.000 141.700 67.400 144.500 ;
        RECT 63.800 141.100 65.800 141.400 ;
        RECT 66.300 141.400 66.600 141.500 ;
        RECT 67.800 141.500 68.200 144.500 ;
        RECT 67.800 141.400 68.100 141.500 ;
        RECT 66.300 141.100 68.100 141.400 ;
        RECT 68.600 141.100 69.000 145.400 ;
        RECT 71.900 145.200 72.200 146.800 ;
        RECT 75.500 146.700 75.900 146.800 ;
        RECT 75.000 146.200 75.400 146.300 ;
        RECT 76.300 146.200 76.700 146.300 ;
        RECT 74.200 145.900 76.700 146.200 ;
        RECT 74.200 145.800 74.600 145.900 ;
        RECT 75.000 145.500 77.800 145.600 ;
        RECT 74.900 145.400 77.800 145.500 ;
        RECT 78.200 145.400 78.600 146.200 ;
        RECT 71.000 144.900 72.200 145.200 ;
        RECT 72.900 145.300 77.800 145.400 ;
        RECT 72.900 145.100 75.300 145.300 ;
        RECT 71.000 144.400 71.300 144.900 ;
        RECT 70.600 144.000 71.300 144.400 ;
        RECT 72.100 144.500 72.500 144.600 ;
        RECT 72.900 144.500 73.200 145.100 ;
        RECT 72.100 144.200 73.200 144.500 ;
        RECT 73.500 144.500 76.200 144.800 ;
        RECT 73.500 144.400 73.900 144.500 ;
        RECT 75.800 144.400 76.200 144.500 ;
        RECT 72.700 143.700 73.100 143.800 ;
        RECT 74.100 143.700 74.500 143.800 ;
        RECT 71.000 143.100 71.400 143.500 ;
        RECT 72.700 143.400 74.500 143.700 ;
        RECT 73.100 143.100 73.400 143.400 ;
        RECT 75.800 143.100 76.200 143.500 ;
        RECT 70.700 141.100 71.300 143.100 ;
        RECT 73.000 141.100 73.400 143.100 ;
        RECT 75.200 142.800 76.200 143.100 ;
        RECT 75.200 141.100 75.600 142.800 ;
        RECT 77.400 141.100 77.800 145.300 ;
        RECT 79.000 145.100 79.300 146.800 ;
        RECT 80.600 145.800 81.000 146.600 ;
        RECT 81.400 145.800 81.800 146.600 ;
        RECT 82.200 146.500 82.900 146.900 ;
        RECT 83.200 146.800 85.000 147.100 ;
        RECT 82.200 145.500 82.500 146.500 ;
        RECT 80.600 145.200 82.500 145.500 ;
        RECT 78.500 144.700 79.400 145.100 ;
        RECT 78.500 141.100 78.900 144.700 ;
        RECT 80.600 143.500 80.900 145.200 ;
        RECT 83.200 144.900 83.500 146.800 ;
        RECT 83.800 146.100 84.200 146.200 ;
        RECT 85.400 146.100 85.800 149.900 ;
        RECT 86.200 148.100 86.600 148.600 ;
        RECT 88.600 148.100 89.000 149.900 ;
        RECT 90.700 149.200 91.300 149.900 ;
        RECT 90.700 148.900 91.400 149.200 ;
        RECT 93.000 148.900 93.400 149.900 ;
        RECT 95.200 149.200 95.600 149.900 ;
        RECT 95.200 148.900 96.200 149.200 ;
        RECT 91.000 148.500 91.400 148.900 ;
        RECT 93.100 148.600 93.400 148.900 ;
        RECT 93.100 148.300 94.500 148.600 ;
        RECT 94.100 148.200 94.500 148.300 ;
        RECT 95.000 148.200 95.400 148.600 ;
        RECT 95.800 148.500 96.200 148.900 ;
        RECT 86.200 147.800 89.000 148.100 ;
        RECT 83.800 145.800 85.800 146.100 ;
        RECT 83.800 145.400 84.200 145.800 ;
        RECT 82.700 144.600 83.500 144.900 ;
        RECT 80.600 141.500 81.000 143.500 ;
        RECT 82.700 141.100 83.100 144.600 ;
        RECT 85.400 141.100 85.800 145.800 ;
        RECT 88.600 147.700 89.000 147.800 ;
        RECT 90.100 147.700 90.500 147.800 ;
        RECT 88.600 147.400 90.500 147.700 ;
        RECT 88.600 145.700 89.000 147.400 ;
        RECT 92.100 147.100 92.500 147.200 ;
        RECT 93.400 147.100 93.800 147.200 ;
        RECT 95.000 147.100 95.300 148.200 ;
        RECT 97.400 147.500 97.800 149.900 ;
        RECT 98.500 148.200 98.900 149.900 ;
        RECT 101.900 149.200 102.700 149.900 ;
        RECT 101.400 148.800 102.700 149.200 ;
        RECT 98.500 147.900 99.400 148.200 ;
        RECT 101.900 147.900 102.700 148.800 ;
        RECT 106.100 147.900 106.900 149.900 ;
        RECT 96.600 147.100 97.400 147.200 ;
        RECT 91.900 146.800 97.400 147.100 ;
        RECT 91.000 146.400 91.400 146.500 ;
        RECT 89.500 146.100 91.400 146.400 ;
        RECT 89.500 146.000 89.900 146.100 ;
        RECT 90.300 145.700 90.700 145.800 ;
        RECT 88.600 145.400 90.700 145.700 ;
        RECT 88.600 141.100 89.000 145.400 ;
        RECT 91.900 145.200 92.200 146.800 ;
        RECT 95.500 146.700 95.900 146.800 ;
        RECT 96.300 146.200 96.700 146.300 ;
        RECT 94.200 145.900 96.700 146.200 ;
        RECT 94.200 145.800 94.600 145.900 ;
        RECT 95.000 145.500 97.800 145.600 ;
        RECT 94.900 145.400 97.800 145.500 ;
        RECT 91.000 144.900 92.200 145.200 ;
        RECT 92.900 145.300 97.800 145.400 ;
        RECT 92.900 145.100 95.300 145.300 ;
        RECT 91.000 144.400 91.300 144.900 ;
        RECT 90.600 144.000 91.300 144.400 ;
        RECT 92.100 144.500 92.500 144.600 ;
        RECT 92.900 144.500 93.200 145.100 ;
        RECT 92.100 144.200 93.200 144.500 ;
        RECT 93.500 144.500 96.200 144.800 ;
        RECT 93.500 144.400 93.900 144.500 ;
        RECT 95.800 144.400 96.200 144.500 ;
        RECT 92.700 143.700 93.100 143.800 ;
        RECT 94.100 143.700 94.500 143.800 ;
        RECT 91.000 143.100 91.400 143.500 ;
        RECT 92.700 143.400 94.500 143.700 ;
        RECT 93.100 143.100 93.400 143.400 ;
        RECT 95.800 143.100 96.200 143.500 ;
        RECT 90.700 141.100 91.300 143.100 ;
        RECT 93.000 141.100 93.400 143.100 ;
        RECT 95.200 142.800 96.200 143.100 ;
        RECT 95.200 141.100 95.600 142.800 ;
        RECT 97.400 141.100 97.800 145.300 ;
        RECT 98.200 144.400 98.600 145.200 ;
        RECT 99.000 141.100 99.400 147.900 ;
        RECT 99.800 146.800 100.200 147.600 ;
        RECT 101.400 146.800 101.800 147.200 ;
        RECT 101.500 146.600 101.800 146.800 ;
        RECT 101.500 146.200 101.900 146.600 ;
        RECT 102.200 146.200 102.500 147.900 ;
        RECT 103.000 147.100 103.400 147.200 ;
        RECT 104.600 147.100 105.000 147.200 ;
        RECT 103.000 146.800 105.000 147.100 ;
        RECT 103.000 146.400 103.400 146.800 ;
        RECT 105.400 146.400 105.800 147.200 ;
        RECT 106.300 146.200 106.600 147.900 ;
        RECT 108.600 147.800 109.000 148.600 ;
        RECT 107.000 146.800 107.400 147.200 ;
        RECT 107.000 146.600 107.300 146.800 ;
        RECT 106.900 146.200 107.300 146.600 ;
        RECT 100.600 145.400 101.000 146.200 ;
        RECT 102.200 145.800 102.600 146.200 ;
        RECT 103.800 146.100 104.200 146.200 ;
        RECT 104.600 146.100 105.000 146.200 ;
        RECT 103.400 145.800 105.400 146.100 ;
        RECT 106.200 145.800 106.600 146.200 ;
        RECT 102.200 145.700 102.500 145.800 ;
        RECT 101.500 145.400 102.500 145.700 ;
        RECT 103.400 145.600 103.800 145.800 ;
        RECT 105.000 145.600 105.400 145.800 ;
        RECT 106.300 145.700 106.600 145.800 ;
        RECT 107.800 146.100 108.200 146.200 ;
        RECT 108.600 146.100 109.000 146.200 ;
        RECT 107.800 145.800 109.000 146.100 ;
        RECT 109.400 146.100 109.800 149.900 ;
        RECT 112.100 149.200 112.500 149.500 ;
        RECT 111.800 148.800 112.500 149.200 ;
        RECT 112.100 148.000 112.500 148.800 ;
        RECT 114.200 148.500 114.600 149.500 ;
        RECT 111.700 147.700 112.500 148.000 ;
        RECT 111.700 147.500 112.100 147.700 ;
        RECT 111.700 147.200 112.000 147.500 ;
        RECT 114.300 147.400 114.600 148.500 ;
        RECT 111.000 146.800 112.000 147.200 ;
        RECT 112.500 147.100 114.600 147.400 ;
        RECT 115.000 148.500 115.400 149.500 ;
        RECT 115.000 147.400 115.300 148.500 ;
        RECT 117.100 148.000 117.500 149.500 ;
        RECT 117.100 147.700 117.900 148.000 ;
        RECT 117.500 147.500 117.900 147.700 ;
        RECT 115.000 147.100 117.100 147.400 ;
        RECT 112.500 146.900 113.000 147.100 ;
        RECT 111.000 146.100 111.400 146.200 ;
        RECT 109.400 145.800 111.400 146.100 ;
        RECT 106.300 145.400 107.300 145.700 ;
        RECT 107.800 145.400 108.200 145.800 ;
        RECT 101.500 145.100 101.800 145.400 ;
        RECT 107.000 145.100 107.300 145.400 ;
        RECT 100.600 141.400 101.000 145.100 ;
        RECT 101.400 141.700 101.800 145.100 ;
        RECT 102.200 144.800 104.200 145.100 ;
        RECT 102.200 141.400 102.600 144.800 ;
        RECT 100.600 141.100 102.600 141.400 ;
        RECT 103.800 141.100 104.200 144.800 ;
        RECT 104.600 144.800 106.600 145.100 ;
        RECT 104.600 141.100 105.000 144.800 ;
        RECT 106.200 141.400 106.600 144.800 ;
        RECT 107.000 141.700 107.400 145.100 ;
        RECT 107.800 141.400 108.200 145.100 ;
        RECT 106.200 141.100 108.200 141.400 ;
        RECT 109.400 141.100 109.800 145.800 ;
        RECT 111.000 145.400 111.400 145.800 ;
        RECT 111.700 144.900 112.000 146.800 ;
        RECT 112.300 146.500 113.000 146.900 ;
        RECT 116.600 146.900 117.100 147.100 ;
        RECT 117.600 147.200 117.900 147.500 ;
        RECT 112.700 145.500 113.000 146.500 ;
        RECT 113.400 145.800 113.800 146.600 ;
        RECT 114.200 145.800 114.600 146.600 ;
        RECT 115.000 145.800 115.400 146.600 ;
        RECT 115.800 145.800 116.200 146.600 ;
        RECT 116.600 146.500 117.300 146.900 ;
        RECT 117.600 146.800 118.600 147.200 ;
        RECT 116.600 145.500 116.900 146.500 ;
        RECT 112.700 145.200 114.600 145.500 ;
        RECT 111.700 144.600 112.500 144.900 ;
        RECT 112.100 141.100 112.500 144.600 ;
        RECT 114.300 143.500 114.600 145.200 ;
        RECT 114.200 141.500 114.600 143.500 ;
        RECT 115.000 145.200 116.900 145.500 ;
        RECT 117.600 145.200 117.900 146.800 ;
        RECT 118.200 146.100 118.600 146.200 ;
        RECT 119.800 146.100 120.200 149.900 ;
        RECT 120.600 148.100 121.000 148.600 ;
        RECT 121.400 148.100 121.800 149.900 ;
        RECT 123.500 149.200 124.100 149.900 ;
        RECT 123.500 148.900 124.200 149.200 ;
        RECT 125.800 148.900 126.200 149.900 ;
        RECT 128.000 149.200 128.400 149.900 ;
        RECT 128.000 148.900 129.000 149.200 ;
        RECT 123.800 148.500 124.200 148.900 ;
        RECT 125.900 148.600 126.200 148.900 ;
        RECT 125.900 148.300 127.300 148.600 ;
        RECT 126.900 148.200 127.300 148.300 ;
        RECT 127.800 148.200 128.200 148.600 ;
        RECT 128.600 148.500 129.000 148.900 ;
        RECT 120.600 147.800 121.800 148.100 ;
        RECT 118.200 145.800 120.200 146.100 ;
        RECT 118.200 145.400 118.600 145.800 ;
        RECT 115.000 143.500 115.300 145.200 ;
        RECT 117.400 144.900 117.900 145.200 ;
        RECT 117.100 144.600 117.900 144.900 ;
        RECT 115.000 141.500 115.400 143.500 ;
        RECT 117.100 141.100 117.500 144.600 ;
        RECT 119.800 141.100 120.200 145.800 ;
        RECT 121.400 147.700 121.800 147.800 ;
        RECT 122.900 147.700 123.300 147.800 ;
        RECT 121.400 147.400 123.300 147.700 ;
        RECT 121.400 145.700 121.800 147.400 ;
        RECT 124.900 147.100 125.300 147.200 ;
        RECT 127.800 147.100 128.100 148.200 ;
        RECT 130.200 147.500 130.600 149.900 ;
        RECT 132.900 148.000 133.300 149.500 ;
        RECT 135.000 148.500 135.400 149.500 ;
        RECT 132.500 147.700 133.300 148.000 ;
        RECT 132.500 147.500 132.900 147.700 ;
        RECT 132.500 147.200 132.800 147.500 ;
        RECT 135.100 147.400 135.400 148.500 ;
        RECT 129.400 147.100 130.200 147.200 ;
        RECT 131.000 147.100 131.400 147.200 ;
        RECT 124.700 146.800 131.400 147.100 ;
        RECT 131.800 146.800 132.800 147.200 ;
        RECT 133.300 147.100 135.400 147.400 ;
        RECT 133.300 146.900 133.800 147.100 ;
        RECT 123.800 146.400 124.200 146.500 ;
        RECT 122.300 146.100 124.200 146.400 ;
        RECT 124.700 146.200 125.000 146.800 ;
        RECT 128.300 146.700 128.700 146.800 ;
        RECT 129.100 146.200 129.500 146.300 ;
        RECT 122.300 146.000 122.700 146.100 ;
        RECT 124.600 145.800 125.000 146.200 ;
        RECT 127.000 145.900 129.500 146.200 ;
        RECT 127.000 145.800 127.400 145.900 ;
        RECT 123.100 145.700 123.500 145.800 ;
        RECT 121.400 145.400 123.500 145.700 ;
        RECT 121.400 141.100 121.800 145.400 ;
        RECT 124.700 145.200 125.000 145.800 ;
        RECT 127.800 145.500 130.600 145.600 ;
        RECT 127.700 145.400 130.600 145.500 ;
        RECT 131.800 145.400 132.200 146.200 ;
        RECT 123.800 144.900 125.000 145.200 ;
        RECT 125.700 145.300 130.600 145.400 ;
        RECT 125.700 145.100 128.100 145.300 ;
        RECT 123.800 144.400 124.100 144.900 ;
        RECT 123.400 144.000 124.100 144.400 ;
        RECT 124.900 144.500 125.300 144.600 ;
        RECT 125.700 144.500 126.000 145.100 ;
        RECT 124.900 144.200 126.000 144.500 ;
        RECT 126.300 144.500 129.000 144.800 ;
        RECT 126.300 144.400 126.700 144.500 ;
        RECT 128.600 144.400 129.000 144.500 ;
        RECT 125.500 143.700 125.900 143.800 ;
        RECT 126.900 143.700 127.300 143.800 ;
        RECT 123.800 143.100 124.200 143.500 ;
        RECT 125.500 143.400 127.300 143.700 ;
        RECT 125.900 143.100 126.200 143.400 ;
        RECT 128.600 143.100 129.000 143.500 ;
        RECT 123.500 141.100 124.100 143.100 ;
        RECT 125.800 141.100 126.200 143.100 ;
        RECT 128.000 142.800 129.000 143.100 ;
        RECT 128.000 141.100 128.400 142.800 ;
        RECT 130.200 141.100 130.600 145.300 ;
        RECT 132.500 145.200 132.800 146.800 ;
        RECT 133.100 146.500 133.800 146.900 ;
        RECT 133.500 145.500 133.800 146.500 ;
        RECT 134.200 145.800 134.600 146.600 ;
        RECT 135.000 145.800 135.400 146.600 ;
        RECT 135.800 146.100 136.200 149.900 ;
        RECT 139.000 149.100 139.400 149.900 ;
        RECT 138.200 148.800 139.400 149.100 ;
        RECT 141.100 149.200 141.700 149.900 ;
        RECT 141.100 148.900 141.800 149.200 ;
        RECT 143.400 148.900 143.800 149.900 ;
        RECT 145.600 149.200 146.000 149.900 ;
        RECT 145.600 148.900 146.600 149.200 ;
        RECT 136.600 148.100 137.000 148.600 ;
        RECT 138.200 148.100 138.500 148.800 ;
        RECT 136.600 147.800 138.500 148.100 ;
        RECT 139.000 147.700 139.400 148.800 ;
        RECT 141.400 148.500 141.800 148.900 ;
        RECT 143.500 148.600 143.800 148.900 ;
        RECT 143.500 148.300 144.900 148.600 ;
        RECT 144.500 148.200 144.900 148.300 ;
        RECT 145.400 148.200 145.800 148.600 ;
        RECT 146.200 148.500 146.600 148.900 ;
        RECT 140.500 147.700 140.900 147.800 ;
        RECT 139.000 147.400 140.900 147.700 ;
        RECT 136.600 146.100 137.000 146.200 ;
        RECT 135.800 145.800 137.000 146.100 ;
        RECT 133.500 145.200 135.400 145.500 ;
        RECT 132.500 144.900 133.000 145.200 ;
        RECT 132.500 144.600 133.300 144.900 ;
        RECT 132.900 141.100 133.300 144.600 ;
        RECT 135.100 143.500 135.400 145.200 ;
        RECT 135.000 141.500 135.400 143.500 ;
        RECT 135.800 141.100 136.200 145.800 ;
        RECT 139.000 145.700 139.400 147.400 ;
        RECT 142.500 147.100 142.900 147.200 ;
        RECT 145.400 147.100 145.700 148.200 ;
        RECT 147.800 147.500 148.200 149.900 ;
        RECT 150.200 147.900 150.600 149.900 ;
        RECT 152.600 148.900 153.000 149.900 ;
        RECT 150.900 148.200 151.300 148.600 ;
        RECT 147.000 147.100 147.800 147.200 ;
        RECT 142.300 146.800 147.800 147.100 ;
        RECT 141.400 146.400 141.800 146.500 ;
        RECT 139.900 146.100 141.800 146.400 ;
        RECT 139.900 146.000 140.300 146.100 ;
        RECT 140.700 145.700 141.100 145.800 ;
        RECT 139.000 145.400 141.100 145.700 ;
        RECT 139.000 141.100 139.400 145.400 ;
        RECT 142.300 145.200 142.600 146.800 ;
        RECT 145.900 146.700 146.300 146.800 ;
        RECT 149.400 146.400 149.800 147.200 ;
        RECT 146.700 146.200 147.100 146.300 ;
        RECT 144.600 145.900 147.100 146.200 ;
        RECT 148.600 146.100 149.000 146.200 ;
        RECT 150.200 146.100 150.500 147.900 ;
        RECT 151.000 147.800 151.400 148.200 ;
        RECT 151.800 147.800 152.200 148.600 ;
        RECT 151.000 147.100 151.300 147.800 ;
        RECT 152.700 147.200 153.000 148.900 ;
        RECT 152.600 147.100 153.000 147.200 ;
        RECT 151.000 146.800 153.000 147.100 ;
        RECT 151.000 146.100 151.400 146.200 ;
        RECT 144.600 145.800 145.000 145.900 ;
        RECT 148.600 145.800 149.400 146.100 ;
        RECT 150.200 145.800 151.400 146.100 ;
        RECT 149.000 145.600 149.400 145.800 ;
        RECT 145.400 145.500 148.200 145.600 ;
        RECT 145.300 145.400 148.200 145.500 ;
        RECT 141.400 144.900 142.600 145.200 ;
        RECT 143.300 145.300 148.200 145.400 ;
        RECT 143.300 145.100 145.700 145.300 ;
        RECT 141.400 144.400 141.700 144.900 ;
        RECT 141.000 144.000 141.700 144.400 ;
        RECT 142.500 144.500 142.900 144.600 ;
        RECT 143.300 144.500 143.600 145.100 ;
        RECT 142.500 144.200 143.600 144.500 ;
        RECT 143.900 144.500 146.600 144.800 ;
        RECT 143.900 144.400 144.300 144.500 ;
        RECT 146.200 144.400 146.600 144.500 ;
        RECT 143.100 143.700 143.500 143.800 ;
        RECT 144.500 143.700 144.900 143.800 ;
        RECT 141.400 143.100 141.800 143.500 ;
        RECT 143.100 143.400 144.900 143.700 ;
        RECT 143.500 143.100 143.800 143.400 ;
        RECT 146.200 143.100 146.600 143.500 ;
        RECT 141.100 141.100 141.700 143.100 ;
        RECT 143.400 141.100 143.800 143.100 ;
        RECT 145.600 142.800 146.600 143.100 ;
        RECT 145.600 141.100 146.000 142.800 ;
        RECT 147.800 141.100 148.200 145.300 ;
        RECT 151.000 145.100 151.300 145.800 ;
        RECT 152.700 145.100 153.000 146.800 ;
        RECT 155.000 148.900 155.400 149.900 ;
        RECT 155.000 147.200 155.300 148.900 ;
        RECT 155.800 147.800 156.200 148.600 ;
        RECT 158.200 147.900 158.600 149.900 ;
        RECT 160.600 148.900 161.000 149.900 ;
        RECT 158.900 148.200 159.300 148.600 ;
        RECT 159.000 148.100 159.400 148.200 ;
        RECT 160.600 148.100 160.900 148.900 ;
        RECT 155.000 146.800 155.400 147.200 ;
        RECT 153.400 146.100 153.800 146.200 ;
        RECT 154.200 146.100 154.600 146.200 ;
        RECT 153.400 145.800 154.600 146.100 ;
        RECT 153.400 145.400 153.800 145.800 ;
        RECT 154.200 145.400 154.600 145.800 ;
        RECT 155.000 145.100 155.300 146.800 ;
        RECT 157.400 146.400 157.800 147.200 ;
        RECT 156.600 146.100 157.000 146.200 ;
        RECT 158.200 146.100 158.500 147.900 ;
        RECT 159.000 147.800 160.900 148.100 ;
        RECT 161.400 147.800 161.800 148.600 ;
        RECT 160.600 147.200 160.900 147.800 ;
        RECT 160.600 146.800 161.000 147.200 ;
        RECT 162.200 146.900 162.600 149.900 ;
        RECT 165.400 148.300 165.800 149.900 ;
        RECT 166.200 148.500 166.600 149.900 ;
        RECT 167.000 148.500 167.400 149.900 ;
        RECT 167.800 148.500 168.200 149.900 ;
        RECT 169.400 148.500 169.800 149.900 ;
        RECT 171.000 148.500 171.400 149.900 ;
        RECT 171.800 148.500 172.200 149.900 ;
        RECT 172.600 148.500 173.000 149.900 ;
        RECT 173.400 148.500 173.800 149.900 ;
        RECT 164.500 147.900 165.800 148.300 ;
        RECT 174.200 148.300 174.600 149.900 ;
        RECT 167.500 147.900 169.800 148.200 ;
        RECT 164.500 147.600 164.900 147.900 ;
        RECT 163.400 147.200 164.900 147.600 ;
        RECT 159.000 146.100 159.400 146.200 ;
        RECT 156.600 145.800 157.400 146.100 ;
        RECT 158.200 145.800 159.400 146.100 ;
        RECT 157.000 145.600 157.400 145.800 ;
        RECT 159.000 145.100 159.300 145.800 ;
        RECT 159.800 145.400 160.200 146.200 ;
        RECT 160.600 145.100 160.900 146.800 ;
        RECT 162.200 146.500 166.600 146.900 ;
        RECT 167.500 146.700 167.900 147.900 ;
        RECT 169.400 147.800 169.800 147.900 ;
        RECT 170.200 147.800 171.000 148.200 ;
        RECT 172.500 147.800 173.000 148.200 ;
        RECT 174.200 147.900 175.400 148.300 ;
        RECT 168.600 146.800 169.000 147.600 ;
        RECT 169.400 147.400 169.800 147.500 ;
        RECT 169.400 147.100 171.600 147.400 ;
        RECT 171.200 147.000 171.600 147.100 ;
        RECT 148.600 144.800 150.600 145.100 ;
        RECT 148.600 141.100 149.000 144.800 ;
        RECT 150.200 141.100 150.600 144.800 ;
        RECT 151.000 141.100 151.400 145.100 ;
        RECT 152.600 144.700 153.500 145.100 ;
        RECT 153.100 141.100 153.500 144.700 ;
        RECT 154.500 144.700 155.400 145.100 ;
        RECT 156.600 144.800 158.600 145.100 ;
        RECT 154.500 142.200 154.900 144.700 ;
        RECT 154.200 141.800 154.900 142.200 ;
        RECT 154.500 141.100 154.900 141.800 ;
        RECT 156.600 141.100 157.000 144.800 ;
        RECT 158.200 141.100 158.600 144.800 ;
        RECT 159.000 141.100 159.400 145.100 ;
        RECT 160.100 144.700 161.000 145.100 ;
        RECT 160.100 141.100 160.500 144.700 ;
        RECT 162.200 143.700 162.600 146.500 ;
        RECT 166.900 146.300 167.900 146.700 ;
        RECT 169.800 146.300 171.400 146.700 ;
        RECT 172.600 146.400 173.000 147.800 ;
        RECT 175.000 147.600 175.400 147.900 ;
        RECT 175.000 147.300 175.900 147.600 ;
        RECT 175.500 146.700 175.900 147.300 ;
        RECT 177.400 147.300 177.800 149.900 ;
        RECT 178.200 148.000 178.600 149.900 ;
        RECT 178.200 147.600 178.700 148.000 ;
        RECT 177.400 147.000 178.000 147.300 ;
        RECT 175.500 146.300 177.400 146.700 ;
        RECT 177.700 146.000 178.000 147.000 ;
        RECT 177.600 145.700 178.000 146.000 ;
        RECT 177.600 144.800 177.900 145.700 ;
        RECT 178.300 145.400 178.700 147.600 ;
        RECT 167.000 144.700 167.400 144.800 ;
        RECT 164.700 144.500 167.400 144.700 ;
        RECT 164.300 144.400 167.400 144.500 ;
        RECT 167.900 144.500 172.200 144.800 ;
        RECT 163.000 144.000 163.800 144.400 ;
        RECT 164.300 144.100 165.000 144.400 ;
        RECT 167.900 144.100 168.200 144.500 ;
        RECT 171.800 144.400 172.200 144.500 ;
        RECT 173.400 144.500 177.900 144.800 ;
        RECT 173.400 144.400 173.800 144.500 ;
        RECT 163.500 143.800 163.800 144.000 ;
        RECT 165.300 143.800 168.200 144.100 ;
        RECT 168.500 143.800 169.800 144.200 ;
        RECT 162.200 143.400 163.200 143.700 ;
        RECT 163.500 143.400 165.600 143.800 ;
        RECT 162.900 143.100 163.200 143.400 ;
        RECT 162.900 142.800 163.400 143.100 ;
        RECT 163.000 141.100 163.400 142.800 ;
        RECT 164.600 141.100 165.000 143.400 ;
        RECT 166.200 141.100 166.600 142.500 ;
        RECT 167.000 141.100 167.400 142.500 ;
        RECT 167.800 141.100 168.200 143.500 ;
        RECT 169.400 141.100 169.800 143.500 ;
        RECT 171.000 141.100 171.400 144.200 ;
        RECT 175.000 143.800 176.300 144.200 ;
        RECT 172.600 143.400 174.700 143.800 ;
        RECT 171.800 141.100 172.200 142.500 ;
        RECT 172.600 141.100 173.000 142.500 ;
        RECT 173.400 141.100 173.800 142.500 ;
        RECT 175.000 141.100 175.400 143.800 ;
        RECT 177.600 143.700 177.900 144.500 ;
        RECT 176.600 143.400 177.900 143.700 ;
        RECT 178.200 145.000 178.700 145.400 ;
        RECT 176.600 141.100 177.000 143.400 ;
        RECT 178.200 141.100 178.600 145.000 ;
        RECT 0.600 135.700 1.000 139.900 ;
        RECT 2.800 138.200 3.200 139.900 ;
        RECT 2.200 137.900 3.200 138.200 ;
        RECT 5.000 137.900 5.400 139.900 ;
        RECT 7.100 137.900 7.700 139.900 ;
        RECT 2.200 137.500 2.600 137.900 ;
        RECT 5.000 137.600 5.300 137.900 ;
        RECT 3.900 137.300 5.700 137.600 ;
        RECT 7.000 137.500 7.400 137.900 ;
        RECT 3.900 137.200 4.300 137.300 ;
        RECT 5.300 137.200 5.700 137.300 ;
        RECT 2.200 136.500 2.600 136.600 ;
        RECT 4.500 136.500 4.900 136.600 ;
        RECT 2.200 136.200 4.900 136.500 ;
        RECT 5.200 136.500 6.300 136.800 ;
        RECT 5.200 135.900 5.500 136.500 ;
        RECT 5.900 136.400 6.300 136.500 ;
        RECT 7.100 136.600 7.800 137.000 ;
        RECT 7.100 136.100 7.400 136.600 ;
        RECT 3.100 135.700 5.500 135.900 ;
        RECT 0.600 135.600 5.500 135.700 ;
        RECT 6.200 135.800 7.400 136.100 ;
        RECT 0.600 135.500 3.500 135.600 ;
        RECT 0.600 135.400 3.400 135.500 ;
        RECT 6.200 135.200 6.500 135.800 ;
        RECT 9.400 135.600 9.800 139.900 ;
        RECT 7.700 135.300 9.800 135.600 ;
        RECT 10.200 135.700 10.600 139.900 ;
        RECT 12.400 138.200 12.800 139.900 ;
        RECT 11.800 137.900 12.800 138.200 ;
        RECT 14.600 137.900 15.000 139.900 ;
        RECT 16.700 137.900 17.300 139.900 ;
        RECT 11.800 137.500 12.200 137.900 ;
        RECT 14.600 137.600 14.900 137.900 ;
        RECT 13.500 137.300 15.300 137.600 ;
        RECT 16.600 137.500 17.000 137.900 ;
        RECT 13.500 137.200 13.900 137.300 ;
        RECT 14.900 137.200 15.300 137.300 ;
        RECT 11.800 136.500 12.200 136.600 ;
        RECT 14.100 136.500 14.500 136.600 ;
        RECT 11.800 136.200 14.500 136.500 ;
        RECT 14.800 136.500 15.900 136.800 ;
        RECT 14.800 135.900 15.100 136.500 ;
        RECT 15.500 136.400 15.900 136.500 ;
        RECT 16.700 136.600 17.400 137.000 ;
        RECT 16.700 136.100 17.000 136.600 ;
        RECT 12.700 135.700 15.100 135.900 ;
        RECT 10.200 135.600 15.100 135.700 ;
        RECT 15.800 135.800 17.000 136.100 ;
        RECT 10.200 135.500 13.100 135.600 ;
        RECT 10.200 135.400 13.000 135.500 ;
        RECT 7.700 135.200 8.100 135.300 ;
        RECT 3.800 135.100 4.200 135.200 ;
        RECT 1.700 134.800 4.200 135.100 ;
        RECT 6.200 134.800 6.600 135.200 ;
        RECT 8.500 134.900 8.900 135.000 ;
        RECT 1.700 134.700 2.100 134.800 ;
        RECT 3.000 134.700 3.400 134.800 ;
        RECT 2.500 134.200 2.900 134.300 ;
        RECT 6.200 134.200 6.500 134.800 ;
        RECT 7.000 134.600 8.900 134.900 ;
        RECT 7.000 134.500 7.400 134.600 ;
        RECT 1.000 133.900 6.500 134.200 ;
        RECT 1.000 133.800 1.800 133.900 ;
        RECT 0.600 131.100 1.000 133.500 ;
        RECT 3.100 132.800 3.400 133.900 ;
        RECT 5.900 133.800 6.300 133.900 ;
        RECT 9.400 133.600 9.800 135.300 ;
        RECT 13.400 135.100 13.800 135.200 ;
        RECT 11.300 134.800 13.800 135.100 ;
        RECT 11.300 134.700 11.700 134.800 ;
        RECT 12.100 134.200 12.500 134.300 ;
        RECT 15.800 134.200 16.100 135.800 ;
        RECT 19.000 135.600 19.400 139.900 ;
        RECT 17.300 135.300 19.400 135.600 ;
        RECT 19.800 137.500 20.200 139.500 ;
        RECT 19.800 135.800 20.100 137.500 ;
        RECT 21.900 136.400 22.300 139.900 ;
        RECT 21.900 136.100 22.700 136.400 ;
        RECT 19.800 135.500 21.700 135.800 ;
        RECT 17.300 135.200 17.700 135.300 ;
        RECT 18.100 134.900 18.500 135.000 ;
        RECT 16.600 134.600 18.500 134.900 ;
        RECT 16.600 134.500 17.000 134.600 ;
        RECT 10.600 133.900 16.200 134.200 ;
        RECT 10.600 133.800 11.400 133.900 ;
        RECT 7.900 133.300 9.800 133.600 ;
        RECT 7.900 133.200 8.300 133.300 ;
        RECT 2.200 132.100 2.600 132.500 ;
        RECT 3.000 132.400 3.400 132.800 ;
        RECT 3.900 132.700 4.300 132.800 ;
        RECT 3.900 132.400 5.300 132.700 ;
        RECT 5.000 132.100 5.300 132.400 ;
        RECT 7.000 132.100 7.400 132.500 ;
        RECT 2.200 131.800 3.200 132.100 ;
        RECT 2.800 131.100 3.200 131.800 ;
        RECT 5.000 131.100 5.400 132.100 ;
        RECT 7.000 131.800 7.700 132.100 ;
        RECT 7.100 131.100 7.700 131.800 ;
        RECT 9.400 131.100 9.800 133.300 ;
        RECT 10.200 131.100 10.600 133.500 ;
        RECT 12.700 132.800 13.000 133.900 ;
        RECT 15.500 133.800 16.200 133.900 ;
        RECT 19.000 133.600 19.400 135.300 ;
        RECT 19.800 134.400 20.200 135.200 ;
        RECT 20.600 134.400 21.000 135.200 ;
        RECT 21.400 134.500 21.700 135.500 ;
        RECT 22.400 135.200 22.700 136.100 ;
        RECT 22.200 134.800 22.700 135.200 ;
        RECT 23.000 135.100 23.400 135.600 ;
        RECT 24.600 135.100 25.000 139.900 ;
        RECT 27.000 137.900 27.400 139.900 ;
        RECT 27.100 137.800 27.400 137.900 ;
        RECT 28.600 137.900 29.000 139.900 ;
        RECT 28.600 137.800 28.900 137.900 ;
        RECT 27.100 137.500 28.900 137.800 ;
        RECT 26.200 137.100 26.600 137.200 ;
        RECT 27.800 137.100 28.200 137.200 ;
        RECT 26.200 136.800 28.200 137.100 ;
        RECT 27.800 136.400 28.200 136.800 ;
        RECT 28.600 136.200 28.900 137.500 ;
        RECT 25.400 136.100 25.800 136.200 ;
        RECT 26.200 136.100 26.600 136.200 ;
        RECT 25.400 135.800 26.600 136.100 ;
        RECT 26.200 135.400 26.600 135.800 ;
        RECT 28.600 135.800 29.000 136.200 ;
        RECT 23.000 134.800 25.000 135.100 ;
        RECT 27.000 134.800 27.800 135.200 ;
        RECT 21.400 134.100 22.100 134.500 ;
        RECT 22.400 134.200 22.700 134.800 ;
        RECT 21.400 133.900 21.900 134.100 ;
        RECT 17.500 133.300 19.400 133.600 ;
        RECT 17.500 133.200 17.900 133.300 ;
        RECT 11.800 132.100 12.200 132.500 ;
        RECT 12.600 132.400 13.000 132.800 ;
        RECT 13.500 132.700 13.900 132.800 ;
        RECT 13.500 132.400 14.900 132.700 ;
        RECT 14.600 132.100 14.900 132.400 ;
        RECT 16.600 132.100 17.000 132.500 ;
        RECT 11.800 131.800 12.800 132.100 ;
        RECT 12.400 131.100 12.800 131.800 ;
        RECT 14.600 131.100 15.000 132.100 ;
        RECT 16.600 131.800 17.300 132.100 ;
        RECT 16.700 131.100 17.300 131.800 ;
        RECT 19.000 131.100 19.400 133.300 ;
        RECT 19.800 133.600 21.900 133.900 ;
        RECT 22.400 133.800 23.400 134.200 ;
        RECT 19.800 132.500 20.100 133.600 ;
        RECT 22.400 133.500 22.700 133.800 ;
        RECT 22.300 133.300 22.700 133.500 ;
        RECT 21.900 133.000 22.700 133.300 ;
        RECT 19.800 131.500 20.200 132.500 ;
        RECT 21.900 131.500 22.300 133.000 ;
        RECT 24.600 131.100 25.000 134.800 ;
        RECT 28.600 134.200 28.900 135.800 ;
        RECT 28.100 134.100 28.900 134.200 ;
        RECT 28.000 133.900 28.900 134.100 ;
        RECT 25.400 132.400 25.800 133.200 ;
        RECT 28.000 131.100 28.400 133.900 ;
        RECT 29.400 133.400 29.800 134.200 ;
        RECT 30.200 134.100 30.600 139.900 ;
        RECT 32.600 137.900 33.000 139.900 ;
        RECT 32.700 137.800 33.000 137.900 ;
        RECT 34.200 137.900 34.600 139.900 ;
        RECT 35.800 137.900 36.200 139.900 ;
        RECT 34.200 137.800 34.500 137.900 ;
        RECT 32.700 137.500 34.500 137.800 ;
        RECT 35.900 137.800 36.200 137.900 ;
        RECT 37.400 137.900 37.800 139.900 ;
        RECT 37.400 137.800 37.700 137.900 ;
        RECT 35.900 137.500 37.700 137.800 ;
        RECT 31.000 135.800 31.400 136.600 ;
        RECT 33.400 136.400 33.800 137.200 ;
        RECT 34.200 136.200 34.500 137.500 ;
        RECT 36.600 136.400 37.000 137.200 ;
        RECT 37.400 136.200 37.700 137.500 ;
        RECT 31.800 135.400 32.200 136.200 ;
        RECT 34.200 136.100 34.600 136.200 ;
        RECT 35.000 136.100 35.400 136.200 ;
        RECT 34.200 135.800 35.400 136.100 ;
        RECT 31.000 134.800 31.400 135.200 ;
        RECT 32.600 134.800 33.400 135.200 ;
        RECT 31.000 134.100 31.300 134.800 ;
        RECT 34.200 134.200 34.500 135.800 ;
        RECT 35.000 135.400 35.400 135.800 ;
        RECT 37.400 135.800 37.800 136.200 ;
        RECT 35.800 134.800 36.600 135.200 ;
        RECT 37.400 134.200 37.700 135.800 ;
        RECT 39.800 135.700 40.200 139.900 ;
        RECT 42.000 138.200 42.400 139.900 ;
        RECT 41.400 137.900 42.400 138.200 ;
        RECT 44.200 137.900 44.600 139.900 ;
        RECT 46.300 137.900 46.900 139.900 ;
        RECT 41.400 137.500 41.800 137.900 ;
        RECT 44.200 137.600 44.500 137.900 ;
        RECT 43.100 137.300 44.900 137.600 ;
        RECT 46.200 137.500 46.600 137.900 ;
        RECT 43.100 137.200 43.500 137.300 ;
        RECT 44.500 137.200 44.900 137.300 ;
        RECT 41.400 136.500 41.800 136.600 ;
        RECT 43.700 136.500 44.100 136.600 ;
        RECT 41.400 136.200 44.100 136.500 ;
        RECT 44.400 136.500 45.500 136.800 ;
        RECT 44.400 135.900 44.700 136.500 ;
        RECT 45.100 136.400 45.500 136.500 ;
        RECT 46.300 136.600 47.000 137.000 ;
        RECT 46.300 136.100 46.600 136.600 ;
        RECT 42.300 135.700 44.700 135.900 ;
        RECT 39.800 135.600 44.700 135.700 ;
        RECT 45.400 135.800 46.600 136.100 ;
        RECT 39.800 135.500 42.700 135.600 ;
        RECT 39.800 135.400 42.600 135.500 ;
        RECT 43.000 135.100 43.400 135.200 ;
        RECT 43.800 135.100 44.200 135.200 ;
        RECT 40.900 134.800 44.200 135.100 ;
        RECT 40.900 134.700 41.300 134.800 ;
        RECT 41.700 134.200 42.100 134.300 ;
        RECT 45.400 134.200 45.700 135.800 ;
        RECT 48.600 135.600 49.000 139.900 ;
        RECT 49.700 136.300 50.100 139.900 ;
        RECT 49.700 135.900 50.600 136.300 ;
        RECT 51.800 135.900 52.200 139.900 ;
        RECT 52.600 136.200 53.000 139.900 ;
        RECT 54.200 136.200 54.600 139.900 ;
        RECT 55.800 137.900 56.200 139.900 ;
        RECT 55.900 137.800 56.200 137.900 ;
        RECT 57.400 137.900 57.800 139.900 ;
        RECT 57.400 137.800 57.700 137.900 ;
        RECT 55.900 137.500 57.700 137.800 ;
        RECT 56.600 136.400 57.000 137.200 ;
        RECT 57.400 136.200 57.700 137.500 ;
        RECT 52.600 135.900 54.600 136.200 ;
        RECT 46.900 135.300 49.000 135.600 ;
        RECT 46.900 135.200 47.300 135.300 ;
        RECT 47.700 134.900 48.100 135.000 ;
        RECT 46.200 134.600 48.100 134.900 ;
        RECT 46.200 134.500 46.600 134.600 ;
        RECT 33.700 134.100 34.500 134.200 ;
        RECT 36.900 134.100 37.700 134.200 ;
        RECT 30.200 133.800 31.300 134.100 ;
        RECT 33.600 133.900 34.500 134.100 ;
        RECT 36.800 133.900 37.700 134.100 ;
        RECT 40.200 133.900 45.700 134.200 ;
        RECT 30.200 133.100 30.600 133.800 ;
        RECT 30.200 132.800 31.100 133.100 ;
        RECT 30.700 131.100 31.100 132.800 ;
        RECT 33.600 131.100 34.000 133.900 ;
        RECT 36.800 133.100 37.200 133.900 ;
        RECT 40.200 133.800 41.000 133.900 ;
        RECT 38.200 133.100 38.600 133.200 ;
        RECT 36.800 132.800 38.600 133.100 ;
        RECT 36.800 131.100 37.200 132.800 ;
        RECT 39.800 131.100 40.200 133.500 ;
        RECT 42.300 132.800 42.600 133.900 ;
        RECT 43.000 133.800 43.400 133.900 ;
        RECT 45.100 133.800 45.500 133.900 ;
        RECT 48.600 133.600 49.000 135.300 ;
        RECT 49.400 134.800 49.800 135.600 ;
        RECT 47.100 133.300 49.000 133.600 ;
        RECT 47.100 133.200 47.500 133.300 ;
        RECT 41.400 132.100 41.800 132.500 ;
        RECT 42.200 132.400 42.600 132.800 ;
        RECT 43.100 132.700 43.500 132.800 ;
        RECT 43.100 132.400 44.500 132.700 ;
        RECT 44.200 132.100 44.500 132.400 ;
        RECT 46.200 132.100 46.600 132.500 ;
        RECT 41.400 131.800 42.400 132.100 ;
        RECT 42.000 131.100 42.400 131.800 ;
        RECT 44.200 131.100 44.600 132.100 ;
        RECT 46.200 131.800 46.900 132.100 ;
        RECT 46.300 131.100 46.900 131.800 ;
        RECT 48.600 131.100 49.000 133.300 ;
        RECT 50.200 134.200 50.500 135.900 ;
        RECT 51.900 135.200 52.200 135.900 ;
        RECT 55.000 135.400 55.400 136.200 ;
        RECT 57.400 135.800 57.800 136.200 ;
        RECT 53.800 135.200 54.200 135.400 ;
        RECT 51.800 134.900 53.000 135.200 ;
        RECT 53.800 134.900 54.600 135.200 ;
        RECT 51.800 134.800 52.200 134.900 ;
        RECT 52.700 134.200 53.000 134.900 ;
        RECT 54.200 134.800 54.600 134.900 ;
        RECT 55.800 134.800 56.600 135.200 ;
        RECT 50.200 134.100 50.600 134.200 ;
        RECT 50.200 133.800 52.100 134.100 ;
        RECT 52.600 133.800 53.000 134.200 ;
        RECT 53.400 133.800 53.800 134.600 ;
        RECT 57.400 134.200 57.700 135.800 ;
        RECT 56.900 134.100 57.700 134.200 ;
        RECT 56.800 133.900 57.700 134.100 ;
        RECT 50.200 132.100 50.500 133.800 ;
        RECT 51.800 133.200 52.100 133.800 ;
        RECT 51.000 132.400 51.400 133.200 ;
        RECT 51.800 132.800 52.200 133.200 ;
        RECT 52.700 133.100 53.000 133.800 ;
        RECT 51.900 132.400 52.300 132.800 ;
        RECT 50.200 131.100 50.600 132.100 ;
        RECT 52.600 131.100 53.000 133.100 ;
        RECT 56.800 131.100 57.200 133.900 ;
        RECT 58.200 133.400 58.600 134.200 ;
        RECT 59.000 133.100 59.400 139.900 ;
        RECT 61.400 137.900 61.800 139.900 ;
        RECT 61.500 137.800 61.800 137.900 ;
        RECT 63.000 137.900 63.400 139.900 ;
        RECT 63.000 137.800 63.300 137.900 ;
        RECT 61.500 137.500 63.300 137.800 ;
        RECT 59.800 135.800 60.200 136.600 ;
        RECT 62.200 136.400 62.600 137.200 ;
        RECT 63.000 136.200 63.300 137.500 ;
        RECT 60.600 135.400 61.000 136.200 ;
        RECT 63.000 135.800 63.400 136.200 ;
        RECT 61.400 134.800 62.200 135.200 ;
        RECT 63.000 134.200 63.300 135.800 ;
        RECT 62.500 134.100 63.300 134.200 ;
        RECT 62.400 133.900 63.300 134.100 ;
        RECT 59.000 132.800 59.900 133.100 ;
        RECT 59.500 132.200 59.900 132.800 ;
        RECT 62.400 132.200 62.800 133.900 ;
        RECT 63.800 133.400 64.200 134.200 ;
        RECT 64.600 133.100 65.000 139.900 ;
        RECT 65.400 135.800 65.800 136.600 ;
        RECT 66.200 135.800 66.600 136.600 ;
        RECT 67.000 133.100 67.400 139.900 ;
        RECT 67.800 133.400 68.200 134.200 ;
        RECT 68.600 133.400 69.000 134.200 ;
        RECT 64.600 132.800 65.500 133.100 ;
        RECT 65.100 132.200 65.500 132.800 ;
        RECT 59.500 131.800 60.200 132.200 ;
        RECT 62.200 131.800 62.800 132.200 ;
        RECT 64.600 131.800 65.500 132.200 ;
        RECT 59.500 131.100 59.900 131.800 ;
        RECT 62.400 131.100 62.800 131.800 ;
        RECT 65.100 131.100 65.500 131.800 ;
        RECT 66.500 132.800 67.400 133.100 ;
        RECT 69.400 133.100 69.800 139.900 ;
        RECT 70.200 135.800 70.600 136.600 ;
        RECT 71.000 136.100 71.400 139.900 ;
        RECT 72.600 137.500 73.000 139.500 ;
        RECT 74.700 139.200 75.100 139.900 ;
        RECT 74.700 138.800 75.400 139.200 ;
        RECT 71.000 135.800 72.100 136.100 ;
        RECT 69.400 132.800 70.300 133.100 ;
        RECT 66.500 132.200 66.900 132.800 ;
        RECT 69.900 132.200 70.300 132.800 ;
        RECT 66.500 131.800 67.400 132.200 ;
        RECT 69.900 131.800 70.600 132.200 ;
        RECT 66.500 131.100 66.900 131.800 ;
        RECT 69.900 131.100 70.300 131.800 ;
        RECT 71.000 131.100 71.400 135.800 ;
        RECT 71.800 135.200 72.100 135.800 ;
        RECT 72.600 135.800 72.900 137.500 ;
        RECT 74.700 136.400 75.100 138.800 ;
        RECT 74.700 136.100 75.500 136.400 ;
        RECT 72.600 135.500 74.500 135.800 ;
        RECT 71.800 134.800 72.200 135.200 ;
        RECT 72.600 134.400 73.000 135.200 ;
        RECT 73.400 134.400 73.800 135.200 ;
        RECT 74.200 134.500 74.500 135.500 ;
        RECT 74.200 134.100 74.900 134.500 ;
        RECT 75.200 134.200 75.500 136.100 ;
        RECT 77.400 135.800 77.800 136.600 ;
        RECT 75.800 134.800 76.200 135.600 ;
        RECT 74.200 133.900 74.700 134.100 ;
        RECT 72.600 133.600 74.700 133.900 ;
        RECT 75.200 133.800 76.200 134.200 ;
        RECT 71.800 132.400 72.200 133.200 ;
        RECT 72.600 132.500 72.900 133.600 ;
        RECT 75.200 133.500 75.500 133.800 ;
        RECT 75.100 133.300 75.500 133.500 ;
        RECT 74.700 133.000 75.500 133.300 ;
        RECT 78.200 133.100 78.600 139.900 ;
        RECT 79.800 135.800 80.200 136.600 ;
        RECT 79.000 133.400 79.400 134.200 ;
        RECT 80.600 133.100 81.000 139.900 ;
        RECT 82.200 136.900 82.600 139.900 ;
        RECT 82.300 136.600 82.600 136.900 ;
        RECT 83.800 139.600 85.800 139.900 ;
        RECT 83.800 136.900 84.200 139.600 ;
        RECT 84.600 136.900 85.000 139.300 ;
        RECT 85.400 137.000 85.800 139.600 ;
        RECT 86.300 139.600 88.100 139.900 ;
        RECT 86.300 139.500 86.600 139.600 ;
        RECT 83.800 136.600 84.100 136.900 ;
        RECT 82.300 136.300 84.100 136.600 ;
        RECT 84.700 136.700 85.000 136.900 ;
        RECT 86.200 136.700 86.600 139.500 ;
        RECT 87.800 139.500 88.100 139.600 ;
        RECT 84.700 136.500 86.600 136.700 ;
        RECT 87.000 136.500 87.400 139.300 ;
        RECT 87.800 136.500 88.200 139.500 ;
        RECT 84.700 136.400 86.500 136.500 ;
        RECT 87.000 136.200 87.300 136.500 ;
        RECT 87.000 136.100 87.400 136.200 ;
        RECT 85.700 135.800 87.400 136.100 ;
        RECT 84.600 134.800 85.400 135.200 ;
        RECT 81.400 133.400 81.800 134.200 ;
        RECT 83.800 133.800 84.600 134.200 ;
        RECT 72.600 131.500 73.000 132.500 ;
        RECT 74.700 131.500 75.100 133.000 ;
        RECT 77.700 132.800 78.600 133.100 ;
        RECT 80.100 132.800 81.000 133.100 ;
        RECT 83.000 132.800 83.900 133.200 ;
        RECT 77.700 132.200 78.100 132.800 ;
        RECT 77.400 131.800 78.100 132.200 ;
        RECT 77.700 131.100 78.100 131.800 ;
        RECT 80.100 132.200 80.500 132.800 ;
        RECT 85.700 132.500 86.000 135.800 ;
        RECT 87.800 135.100 88.200 135.200 ;
        RECT 91.000 135.100 91.400 139.900 ;
        RECT 91.800 135.800 92.200 136.600 ;
        RECT 92.600 136.200 93.000 139.900 ;
        RECT 94.200 139.600 96.200 139.900 ;
        RECT 94.200 136.200 94.600 139.600 ;
        RECT 92.600 135.900 94.600 136.200 ;
        RECT 95.000 135.900 95.400 139.300 ;
        RECT 95.800 135.900 96.200 139.600 ;
        RECT 95.000 135.600 95.300 135.900 ;
        RECT 96.600 135.600 97.000 139.900 ;
        RECT 98.700 137.900 99.300 139.900 ;
        RECT 101.000 137.900 101.400 139.900 ;
        RECT 103.200 138.200 103.600 139.900 ;
        RECT 103.200 137.900 104.200 138.200 ;
        RECT 99.000 137.500 99.400 137.900 ;
        RECT 101.100 137.600 101.400 137.900 ;
        RECT 100.700 137.300 102.500 137.600 ;
        RECT 103.800 137.500 104.200 137.900 ;
        RECT 100.700 137.200 101.100 137.300 ;
        RECT 102.100 137.200 102.500 137.300 ;
        RECT 98.600 136.600 99.300 137.000 ;
        RECT 99.000 136.100 99.300 136.600 ;
        RECT 100.100 136.500 101.200 136.800 ;
        RECT 100.100 136.400 100.500 136.500 ;
        RECT 99.000 135.800 100.200 136.100 ;
        RECT 93.000 135.200 93.400 135.400 ;
        RECT 94.300 135.300 95.300 135.600 ;
        RECT 94.300 135.200 94.600 135.300 ;
        RECT 87.800 134.800 91.400 135.100 ;
        RECT 92.600 134.900 93.400 135.200 ;
        RECT 92.600 134.800 93.000 134.900 ;
        RECT 94.200 134.800 94.600 135.200 ;
        RECT 95.800 134.800 96.200 135.600 ;
        RECT 96.600 135.300 98.700 135.600 ;
        RECT 87.800 134.100 88.200 134.200 ;
        RECT 90.200 134.100 90.600 134.200 ;
        RECT 87.800 133.800 90.600 134.100 ;
        RECT 90.200 133.400 90.600 133.800 ;
        RECT 91.000 133.100 91.400 134.800 ;
        RECT 93.400 133.800 93.800 134.600 ;
        RECT 94.300 133.100 94.600 134.800 ;
        RECT 94.900 134.400 95.300 134.800 ;
        RECT 95.000 134.200 95.300 134.400 ;
        RECT 95.000 133.800 95.400 134.200 ;
        RECT 96.600 133.600 97.000 135.300 ;
        RECT 98.300 135.200 98.700 135.300 ;
        RECT 97.500 134.900 97.900 135.000 ;
        RECT 97.500 134.600 99.400 134.900 ;
        RECT 99.000 134.500 99.400 134.600 ;
        RECT 99.900 134.200 100.200 135.800 ;
        RECT 100.900 135.900 101.200 136.500 ;
        RECT 101.500 136.500 101.900 136.600 ;
        RECT 103.800 136.500 104.200 136.600 ;
        RECT 101.500 136.200 104.200 136.500 ;
        RECT 100.900 135.700 103.300 135.900 ;
        RECT 105.400 135.700 105.800 139.900 ;
        RECT 106.200 136.200 106.600 139.900 ;
        RECT 107.800 139.600 109.800 139.900 ;
        RECT 107.800 136.200 108.200 139.600 ;
        RECT 106.200 135.900 108.200 136.200 ;
        RECT 108.600 135.900 109.000 139.300 ;
        RECT 109.400 135.900 109.800 139.600 ;
        RECT 100.900 135.600 105.800 135.700 ;
        RECT 108.600 135.600 108.900 135.900 ;
        RECT 102.900 135.500 105.800 135.600 ;
        RECT 103.000 135.400 105.800 135.500 ;
        RECT 106.600 135.200 107.000 135.400 ;
        RECT 107.900 135.300 108.900 135.600 ;
        RECT 107.900 135.200 108.200 135.300 ;
        RECT 102.200 135.100 102.600 135.200 ;
        RECT 102.200 134.800 104.700 135.100 ;
        RECT 106.200 134.900 107.000 135.200 ;
        RECT 106.200 134.800 106.600 134.900 ;
        RECT 107.800 134.800 108.200 135.200 ;
        RECT 109.400 135.100 109.800 135.600 ;
        RECT 110.200 135.100 110.600 135.200 ;
        RECT 109.400 134.800 110.600 135.100 ;
        RECT 111.000 135.100 111.400 139.900 ;
        RECT 113.700 136.400 114.100 139.900 ;
        RECT 115.800 137.500 116.200 139.500 ;
        RECT 113.300 136.100 114.100 136.400 ;
        RECT 112.600 135.100 113.000 135.600 ;
        RECT 111.000 134.800 113.000 135.100 ;
        RECT 103.000 134.700 103.400 134.800 ;
        RECT 104.300 134.700 104.700 134.800 ;
        RECT 103.500 134.200 103.900 134.300 ;
        RECT 99.900 133.900 105.400 134.200 ;
        RECT 100.100 133.800 100.500 133.900 ;
        RECT 103.000 133.800 103.400 133.900 ;
        RECT 104.600 133.800 105.400 133.900 ;
        RECT 107.000 133.800 107.400 134.600 ;
        RECT 96.600 133.300 98.500 133.600 ;
        RECT 91.000 132.800 91.900 133.100 ;
        RECT 84.000 132.200 86.000 132.500 ;
        RECT 80.100 131.800 81.000 132.200 ;
        RECT 84.000 132.100 84.300 132.200 ;
        RECT 83.800 131.800 84.300 132.100 ;
        RECT 85.400 132.100 86.000 132.200 ;
        RECT 88.600 132.100 89.000 132.200 ;
        RECT 85.400 131.800 89.000 132.100 ;
        RECT 80.100 131.100 80.500 131.800 ;
        RECT 83.800 131.100 84.200 131.800 ;
        RECT 85.400 131.100 85.800 131.800 ;
        RECT 91.500 131.100 91.900 132.800 ;
        RECT 94.100 131.100 94.900 133.100 ;
        RECT 96.600 131.100 97.000 133.300 ;
        RECT 98.100 133.200 98.500 133.300 ;
        RECT 103.000 132.800 103.300 133.800 ;
        RECT 102.100 132.700 102.500 132.800 ;
        RECT 99.000 132.100 99.400 132.500 ;
        RECT 101.100 132.400 102.500 132.700 ;
        RECT 103.000 132.400 103.400 132.800 ;
        RECT 101.100 132.100 101.400 132.400 ;
        RECT 103.800 132.100 104.200 132.500 ;
        RECT 98.700 131.800 99.400 132.100 ;
        RECT 98.700 131.100 99.300 131.800 ;
        RECT 101.000 131.100 101.400 132.100 ;
        RECT 103.200 131.800 104.200 132.100 ;
        RECT 103.200 131.100 103.600 131.800 ;
        RECT 105.400 131.100 105.800 133.500 ;
        RECT 107.900 133.100 108.200 134.800 ;
        RECT 108.500 134.400 108.900 134.800 ;
        RECT 108.600 134.200 108.900 134.400 ;
        RECT 108.600 133.800 109.000 134.200 ;
        RECT 107.700 131.100 108.500 133.100 ;
        RECT 110.200 132.400 110.600 133.200 ;
        RECT 111.000 131.100 111.400 134.800 ;
        RECT 113.300 134.200 113.600 136.100 ;
        RECT 115.900 135.800 116.200 137.500 ;
        RECT 114.300 135.500 116.200 135.800 ;
        RECT 116.600 135.700 117.000 139.900 ;
        RECT 118.800 138.200 119.200 139.900 ;
        RECT 118.200 137.900 119.200 138.200 ;
        RECT 121.000 137.900 121.400 139.900 ;
        RECT 123.100 137.900 123.700 139.900 ;
        RECT 118.200 137.500 118.600 137.900 ;
        RECT 121.000 137.600 121.300 137.900 ;
        RECT 119.900 137.300 121.700 137.600 ;
        RECT 123.000 137.500 123.400 137.900 ;
        RECT 119.900 137.200 120.300 137.300 ;
        RECT 121.300 137.200 121.700 137.300 ;
        RECT 118.200 136.500 118.600 136.600 ;
        RECT 120.500 136.500 120.900 136.600 ;
        RECT 118.200 136.200 120.900 136.500 ;
        RECT 121.200 136.500 122.300 136.800 ;
        RECT 121.200 135.900 121.500 136.500 ;
        RECT 121.900 136.400 122.300 136.500 ;
        RECT 123.100 136.600 123.800 137.000 ;
        RECT 123.100 136.100 123.400 136.600 ;
        RECT 119.100 135.700 121.500 135.900 ;
        RECT 116.600 135.600 121.500 135.700 ;
        RECT 122.200 135.800 123.400 136.100 ;
        RECT 116.600 135.500 119.500 135.600 ;
        RECT 114.300 134.500 114.600 135.500 ;
        RECT 116.600 135.400 119.400 135.500 ;
        RECT 112.600 133.800 113.600 134.200 ;
        RECT 113.900 134.100 114.600 134.500 ;
        RECT 115.000 134.400 115.400 135.200 ;
        RECT 115.800 134.400 116.200 135.200 ;
        RECT 119.800 135.100 120.200 135.200 ;
        RECT 117.700 134.800 120.200 135.100 ;
        RECT 117.700 134.700 118.100 134.800 ;
        RECT 118.500 134.200 118.900 134.300 ;
        RECT 122.200 134.200 122.500 135.800 ;
        RECT 125.400 135.600 125.800 139.900 ;
        RECT 123.700 135.300 125.800 135.600 ;
        RECT 123.700 135.200 124.100 135.300 ;
        RECT 124.500 134.900 124.900 135.000 ;
        RECT 123.000 134.600 124.900 134.900 ;
        RECT 123.000 134.500 123.400 134.600 ;
        RECT 113.300 133.500 113.600 133.800 ;
        RECT 114.100 133.900 114.600 134.100 ;
        RECT 117.000 133.900 122.500 134.200 ;
        RECT 114.100 133.600 116.200 133.900 ;
        RECT 117.000 133.800 117.800 133.900 ;
        RECT 119.000 133.800 119.400 133.900 ;
        RECT 121.900 133.800 122.300 133.900 ;
        RECT 113.300 133.300 113.700 133.500 ;
        RECT 113.300 133.000 114.100 133.300 ;
        RECT 113.700 132.200 114.100 133.000 ;
        RECT 115.900 132.500 116.200 133.600 ;
        RECT 113.400 131.800 114.100 132.200 ;
        RECT 113.700 131.500 114.100 131.800 ;
        RECT 115.800 131.500 116.200 132.500 ;
        RECT 116.600 131.100 117.000 133.500 ;
        RECT 119.100 132.800 119.400 133.800 ;
        RECT 125.400 133.600 125.800 135.300 ;
        RECT 126.200 135.100 126.600 135.200 ;
        RECT 127.000 135.100 127.400 139.900 ;
        RECT 129.700 136.400 130.100 139.900 ;
        RECT 131.800 137.500 132.200 139.500 ;
        RECT 129.300 136.100 130.100 136.400 ;
        RECT 126.200 134.800 127.400 135.100 ;
        RECT 127.800 135.100 128.200 135.200 ;
        RECT 128.600 135.100 129.000 135.600 ;
        RECT 127.800 134.800 129.000 135.100 ;
        RECT 123.900 133.300 125.800 133.600 ;
        RECT 123.900 133.200 124.300 133.300 ;
        RECT 125.400 133.100 125.800 133.300 ;
        RECT 126.200 133.100 126.600 133.200 ;
        RECT 125.400 132.800 126.600 133.100 ;
        RECT 118.200 132.100 118.600 132.500 ;
        RECT 119.000 132.400 119.400 132.800 ;
        RECT 119.900 132.700 120.300 132.800 ;
        RECT 119.900 132.400 121.300 132.700 ;
        RECT 121.000 132.100 121.300 132.400 ;
        RECT 123.000 132.100 123.400 132.500 ;
        RECT 118.200 131.800 119.200 132.100 ;
        RECT 118.800 131.100 119.200 131.800 ;
        RECT 121.000 131.100 121.400 132.100 ;
        RECT 123.000 131.800 123.700 132.100 ;
        RECT 123.100 131.100 123.700 131.800 ;
        RECT 125.400 131.100 125.800 132.800 ;
        RECT 126.200 132.400 126.600 132.800 ;
        RECT 127.000 131.100 127.400 134.800 ;
        RECT 129.300 134.200 129.600 136.100 ;
        RECT 131.900 135.800 132.200 137.500 ;
        RECT 134.500 136.400 134.900 139.900 ;
        RECT 136.600 137.500 137.000 139.500 ;
        RECT 130.300 135.500 132.200 135.800 ;
        RECT 134.100 136.100 134.900 136.400 ;
        RECT 130.300 134.500 130.600 135.500 ;
        RECT 127.800 134.100 128.200 134.200 ;
        RECT 128.600 134.100 129.600 134.200 ;
        RECT 129.900 134.100 130.600 134.500 ;
        RECT 131.000 134.400 131.400 135.200 ;
        RECT 131.800 134.400 132.200 135.200 ;
        RECT 132.600 135.100 133.000 135.200 ;
        RECT 133.400 135.100 133.800 135.600 ;
        RECT 132.600 134.800 133.800 135.100 ;
        RECT 134.100 135.200 134.400 136.100 ;
        RECT 136.700 135.800 137.000 137.500 ;
        RECT 135.100 135.500 137.000 135.800 ;
        RECT 139.000 135.600 139.400 139.900 ;
        RECT 141.100 137.900 141.700 139.900 ;
        RECT 143.400 137.900 143.800 139.900 ;
        RECT 145.600 138.200 146.000 139.900 ;
        RECT 145.600 137.900 146.600 138.200 ;
        RECT 141.400 137.500 141.800 137.900 ;
        RECT 143.500 137.600 143.800 137.900 ;
        RECT 143.100 137.300 144.900 137.600 ;
        RECT 146.200 137.500 146.600 137.900 ;
        RECT 143.100 137.200 143.500 137.300 ;
        RECT 144.500 137.200 144.900 137.300 ;
        RECT 141.000 136.600 141.700 137.000 ;
        RECT 141.400 136.100 141.700 136.600 ;
        RECT 142.500 136.500 143.600 136.800 ;
        RECT 142.500 136.400 142.900 136.500 ;
        RECT 141.400 135.800 142.600 136.100 ;
        RECT 134.100 134.800 134.600 135.200 ;
        RECT 134.100 134.200 134.400 134.800 ;
        RECT 135.100 134.500 135.400 135.500 ;
        RECT 139.000 135.300 141.100 135.600 ;
        RECT 127.800 133.800 129.600 134.100 ;
        RECT 129.300 133.500 129.600 133.800 ;
        RECT 130.100 133.900 130.600 134.100 ;
        RECT 130.100 133.600 132.200 133.900 ;
        RECT 133.400 133.800 134.400 134.200 ;
        RECT 134.700 134.100 135.400 134.500 ;
        RECT 135.800 134.400 136.200 135.200 ;
        RECT 136.600 135.100 137.000 135.200 ;
        RECT 137.400 135.100 137.800 135.200 ;
        RECT 136.600 134.800 137.800 135.100 ;
        RECT 136.600 134.400 137.000 134.800 ;
        RECT 129.300 133.300 129.700 133.500 ;
        RECT 129.300 133.000 130.100 133.300 ;
        RECT 129.700 131.500 130.100 133.000 ;
        RECT 131.900 132.500 132.200 133.600 ;
        RECT 134.100 133.500 134.400 133.800 ;
        RECT 134.900 133.900 135.400 134.100 ;
        RECT 134.900 133.600 137.000 133.900 ;
        RECT 134.100 133.300 134.500 133.500 ;
        RECT 134.100 133.000 134.900 133.300 ;
        RECT 131.800 131.500 132.200 132.500 ;
        RECT 134.500 131.500 134.900 133.000 ;
        RECT 136.700 132.500 137.000 133.600 ;
        RECT 136.600 131.500 137.000 132.500 ;
        RECT 139.000 133.600 139.400 135.300 ;
        RECT 140.700 135.200 141.100 135.300 ;
        RECT 139.900 134.900 140.300 135.000 ;
        RECT 139.900 134.600 141.800 134.900 ;
        RECT 141.400 134.500 141.800 134.600 ;
        RECT 142.300 134.200 142.600 135.800 ;
        RECT 143.300 135.900 143.600 136.500 ;
        RECT 143.900 136.500 144.300 136.600 ;
        RECT 146.200 136.500 146.600 136.600 ;
        RECT 143.900 136.200 146.600 136.500 ;
        RECT 143.300 135.700 145.700 135.900 ;
        RECT 147.800 135.700 148.200 139.900 ;
        RECT 149.000 136.800 149.400 137.200 ;
        RECT 149.000 136.200 149.300 136.800 ;
        RECT 149.700 136.200 150.100 139.900 ;
        RECT 148.600 135.900 149.300 136.200 ;
        RECT 149.600 135.900 150.100 136.200 ;
        RECT 148.600 135.800 149.000 135.900 ;
        RECT 143.300 135.600 148.200 135.700 ;
        RECT 145.300 135.500 148.200 135.600 ;
        RECT 145.400 135.400 148.200 135.500 ;
        RECT 144.600 135.100 145.000 135.200 ;
        RECT 144.600 134.800 147.100 135.100 ;
        RECT 146.700 134.700 147.100 134.800 ;
        RECT 145.900 134.200 146.300 134.300 ;
        RECT 149.600 134.200 149.900 135.900 ;
        RECT 150.200 135.100 150.600 135.200 ;
        RECT 152.600 135.100 153.000 139.900 ;
        RECT 155.300 136.400 155.700 139.900 ;
        RECT 157.400 137.500 157.800 139.500 ;
        RECT 154.900 136.100 155.700 136.400 ;
        RECT 154.200 135.100 154.600 135.600 ;
        RECT 150.200 134.800 154.600 135.100 ;
        RECT 150.200 134.400 150.600 134.800 ;
        RECT 142.300 133.900 147.800 134.200 ;
        RECT 142.500 133.800 142.900 133.900 ;
        RECT 139.000 133.300 140.900 133.600 ;
        RECT 139.000 131.100 139.400 133.300 ;
        RECT 140.500 133.200 140.900 133.300 ;
        RECT 145.400 132.800 145.700 133.900 ;
        RECT 147.000 133.800 147.800 133.900 ;
        RECT 148.600 133.800 149.900 134.200 ;
        RECT 151.000 134.100 151.400 134.200 ;
        RECT 150.600 133.800 151.400 134.100 ;
        RECT 144.500 132.700 144.900 132.800 ;
        RECT 141.400 132.100 141.800 132.500 ;
        RECT 143.500 132.400 144.900 132.700 ;
        RECT 145.400 132.400 145.800 132.800 ;
        RECT 143.500 132.100 143.800 132.400 ;
        RECT 146.200 132.100 146.600 132.500 ;
        RECT 141.100 131.800 141.800 132.100 ;
        RECT 141.100 131.100 141.700 131.800 ;
        RECT 143.400 131.100 143.800 132.100 ;
        RECT 145.600 131.800 146.600 132.100 ;
        RECT 145.600 131.100 146.000 131.800 ;
        RECT 147.800 131.100 148.200 133.500 ;
        RECT 148.700 133.100 149.000 133.800 ;
        RECT 150.600 133.600 151.000 133.800 ;
        RECT 149.500 133.100 151.300 133.300 ;
        RECT 148.600 131.100 149.000 133.100 ;
        RECT 149.400 133.000 151.400 133.100 ;
        RECT 149.400 131.100 149.800 133.000 ;
        RECT 151.000 131.100 151.400 133.000 ;
        RECT 151.800 132.400 152.200 133.200 ;
        RECT 152.600 131.100 153.000 134.800 ;
        RECT 154.900 134.200 155.200 136.100 ;
        RECT 157.500 135.800 157.800 137.500 ;
        RECT 158.200 136.900 158.600 139.900 ;
        RECT 158.300 136.600 158.600 136.900 ;
        RECT 159.800 139.600 161.800 139.900 ;
        RECT 159.800 136.900 160.200 139.600 ;
        RECT 160.600 136.900 161.000 139.300 ;
        RECT 161.400 137.000 161.800 139.600 ;
        RECT 162.300 139.600 164.100 139.900 ;
        RECT 162.300 139.500 162.600 139.600 ;
        RECT 159.800 136.600 160.100 136.900 ;
        RECT 158.300 136.300 160.100 136.600 ;
        RECT 160.700 136.700 161.000 136.900 ;
        RECT 162.200 136.700 162.600 139.500 ;
        RECT 163.800 139.500 164.100 139.600 ;
        RECT 160.700 136.500 162.600 136.700 ;
        RECT 163.000 136.500 163.400 139.300 ;
        RECT 163.800 136.500 164.200 139.500 ;
        RECT 165.000 136.800 165.400 137.200 ;
        RECT 160.700 136.400 162.500 136.500 ;
        RECT 163.000 136.200 163.300 136.500 ;
        RECT 165.000 136.200 165.300 136.800 ;
        RECT 165.700 136.200 166.100 139.900 ;
        RECT 163.000 136.100 163.400 136.200 ;
        RECT 155.900 135.500 157.800 135.800 ;
        RECT 161.700 135.800 163.400 136.100 ;
        RECT 163.800 136.100 164.200 136.200 ;
        RECT 164.600 136.100 165.300 136.200 ;
        RECT 163.800 135.900 165.300 136.100 ;
        RECT 165.600 135.900 166.100 136.200 ;
        RECT 167.800 137.500 168.200 139.500 ;
        RECT 163.800 135.800 165.000 135.900 ;
        RECT 155.900 134.500 156.200 135.500 ;
        RECT 154.200 133.800 155.200 134.200 ;
        RECT 155.500 134.100 156.200 134.500 ;
        RECT 156.600 134.400 157.000 135.200 ;
        RECT 157.400 134.400 157.800 135.200 ;
        RECT 160.600 134.800 161.400 135.200 ;
        RECT 154.900 133.500 155.200 133.800 ;
        RECT 155.700 133.900 156.200 134.100 ;
        RECT 155.700 133.600 157.800 133.900 ;
        RECT 159.800 133.800 160.600 134.200 ;
        RECT 154.900 133.300 155.300 133.500 ;
        RECT 154.900 133.000 155.700 133.300 ;
        RECT 155.300 132.200 155.700 133.000 ;
        RECT 157.500 132.500 157.800 133.600 ;
        RECT 159.000 132.800 160.200 133.200 ;
        RECT 161.700 132.500 162.000 135.800 ;
        RECT 163.000 135.100 163.400 135.200 ;
        RECT 165.600 135.100 165.900 135.900 ;
        RECT 167.800 135.800 168.100 137.500 ;
        RECT 169.900 136.400 170.300 139.900 ;
        RECT 172.600 137.500 173.000 139.500 ;
        RECT 174.700 139.200 175.100 139.900 ;
        RECT 174.200 138.800 175.100 139.200 ;
        RECT 169.900 136.100 170.700 136.400 ;
        RECT 167.800 135.500 169.700 135.800 ;
        RECT 163.000 134.800 165.900 135.100 ;
        RECT 165.600 134.200 165.900 134.800 ;
        RECT 166.200 134.400 166.600 135.200 ;
        RECT 167.800 134.400 168.200 135.200 ;
        RECT 168.600 134.400 169.000 135.200 ;
        RECT 169.400 134.500 169.700 135.500 ;
        RECT 164.600 133.800 165.900 134.200 ;
        RECT 167.000 134.100 167.400 134.200 ;
        RECT 166.600 133.800 167.400 134.100 ;
        RECT 169.400 134.100 170.100 134.500 ;
        RECT 170.400 134.200 170.700 136.100 ;
        RECT 172.600 135.800 172.900 137.500 ;
        RECT 174.700 136.400 175.100 138.800 ;
        RECT 174.700 136.100 175.500 136.400 ;
        RECT 171.000 134.800 171.400 135.600 ;
        RECT 172.600 135.500 174.500 135.800 ;
        RECT 172.600 134.400 173.000 135.200 ;
        RECT 173.400 134.400 173.800 135.200 ;
        RECT 174.200 134.500 174.500 135.500 ;
        RECT 169.400 133.900 169.900 134.100 ;
        RECT 164.700 133.100 165.000 133.800 ;
        RECT 166.600 133.600 167.000 133.800 ;
        RECT 167.800 133.600 169.900 133.900 ;
        RECT 170.400 133.800 171.400 134.200 ;
        RECT 174.200 134.100 174.900 134.500 ;
        RECT 175.200 134.200 175.500 136.100 ;
        RECT 175.800 135.100 176.200 135.600 ;
        RECT 177.400 135.100 177.800 139.900 ;
        RECT 175.800 134.800 177.800 135.100 ;
        RECT 178.200 135.800 178.600 136.200 ;
        RECT 178.200 135.100 178.500 135.800 ;
        RECT 179.000 135.100 179.400 139.900 ;
        RECT 178.200 134.800 179.400 135.100 ;
        RECT 174.200 133.900 174.700 134.100 ;
        RECT 165.500 133.100 167.300 133.300 ;
        RECT 155.000 131.800 155.700 132.200 ;
        RECT 155.300 131.500 155.700 131.800 ;
        RECT 157.400 131.500 157.800 132.500 ;
        RECT 160.000 132.200 162.000 132.500 ;
        RECT 160.000 132.100 160.300 132.200 ;
        RECT 159.800 131.800 160.300 132.100 ;
        RECT 161.400 132.100 162.000 132.200 ;
        RECT 159.800 131.100 160.200 131.800 ;
        RECT 161.400 131.100 161.800 132.100 ;
        RECT 164.600 131.100 165.000 133.100 ;
        RECT 165.400 133.000 167.400 133.100 ;
        RECT 165.400 131.100 165.800 133.000 ;
        RECT 167.000 131.100 167.400 133.000 ;
        RECT 167.800 132.500 168.100 133.600 ;
        RECT 170.400 133.500 170.700 133.800 ;
        RECT 170.300 133.300 170.700 133.500 ;
        RECT 169.900 133.000 170.700 133.300 ;
        RECT 172.600 133.600 174.700 133.900 ;
        RECT 175.200 133.800 176.200 134.200 ;
        RECT 167.800 131.500 168.200 132.500 ;
        RECT 169.900 132.200 170.300 133.000 ;
        RECT 169.400 131.800 170.300 132.200 ;
        RECT 169.900 131.500 170.300 131.800 ;
        RECT 172.600 132.500 172.900 133.600 ;
        RECT 175.200 133.500 175.500 133.800 ;
        RECT 175.100 133.300 175.500 133.500 ;
        RECT 174.700 133.000 175.500 133.300 ;
        RECT 172.600 131.500 173.000 132.500 ;
        RECT 174.700 131.500 175.100 133.000 ;
        RECT 177.400 131.100 177.800 134.800 ;
        RECT 178.200 133.800 178.600 134.200 ;
        RECT 178.200 133.200 178.500 133.800 ;
        RECT 178.200 132.400 178.600 133.200 ;
        RECT 179.000 131.100 179.400 134.800 ;
        RECT 179.800 132.400 180.200 133.200 ;
        RECT 2.500 129.200 2.900 129.500 ;
        RECT 2.500 128.800 3.400 129.200 ;
        RECT 2.500 128.000 2.900 128.800 ;
        RECT 4.600 128.500 5.000 129.500 ;
        RECT 2.100 127.700 2.900 128.000 ;
        RECT 2.100 127.500 2.500 127.700 ;
        RECT 2.100 127.200 2.400 127.500 ;
        RECT 4.700 127.400 5.000 128.500 ;
        RECT 1.400 126.800 2.400 127.200 ;
        RECT 2.900 127.100 5.000 127.400 ;
        RECT 2.900 126.900 3.400 127.100 ;
        RECT 1.400 125.400 1.800 126.200 ;
        RECT 2.100 124.900 2.400 126.800 ;
        RECT 2.700 126.500 3.400 126.900 ;
        RECT 3.100 125.500 3.400 126.500 ;
        RECT 3.800 125.800 4.200 126.600 ;
        RECT 4.600 125.800 5.000 126.600 ;
        RECT 5.400 126.100 5.800 129.900 ;
        RECT 6.200 127.800 6.600 128.600 ;
        RECT 7.000 128.500 7.400 129.500 ;
        RECT 7.000 127.400 7.300 128.500 ;
        RECT 9.100 128.000 9.500 129.500 ;
        RECT 9.100 127.700 9.900 128.000 ;
        RECT 9.500 127.500 9.900 127.700 ;
        RECT 7.000 127.100 9.100 127.400 ;
        RECT 8.600 126.900 9.100 127.100 ;
        RECT 9.600 127.200 9.900 127.500 ;
        RECT 9.600 127.100 10.600 127.200 ;
        RECT 11.000 127.100 11.400 127.200 ;
        RECT 6.200 126.100 6.600 126.200 ;
        RECT 5.400 125.800 6.600 126.100 ;
        RECT 7.000 125.800 7.400 126.600 ;
        RECT 7.800 125.800 8.200 126.600 ;
        RECT 8.600 126.500 9.300 126.900 ;
        RECT 9.600 126.800 11.400 127.100 ;
        RECT 3.100 125.200 5.000 125.500 ;
        RECT 2.100 124.600 2.900 124.900 ;
        RECT 2.500 121.100 2.900 124.600 ;
        RECT 4.700 123.500 5.000 125.200 ;
        RECT 4.600 121.500 5.000 123.500 ;
        RECT 5.400 121.100 5.800 125.800 ;
        RECT 8.600 125.500 8.900 126.500 ;
        RECT 7.000 125.200 8.900 125.500 ;
        RECT 7.000 123.500 7.300 125.200 ;
        RECT 9.600 124.900 9.900 126.800 ;
        RECT 10.200 126.100 10.600 126.200 ;
        RECT 11.800 126.100 12.200 129.900 ;
        RECT 12.600 127.800 13.000 128.600 ;
        RECT 13.400 127.500 13.800 129.900 ;
        RECT 15.600 129.200 16.000 129.900 ;
        RECT 15.000 128.900 16.000 129.200 ;
        RECT 17.800 128.900 18.200 129.900 ;
        RECT 19.900 129.200 20.500 129.900 ;
        RECT 19.800 128.900 20.500 129.200 ;
        RECT 15.000 128.500 15.400 128.900 ;
        RECT 17.800 128.600 18.100 128.900 ;
        RECT 15.800 127.800 16.200 128.600 ;
        RECT 16.700 128.300 18.100 128.600 ;
        RECT 19.800 128.500 20.200 128.900 ;
        RECT 16.700 128.200 17.100 128.300 ;
        RECT 12.600 127.100 13.000 127.200 ;
        RECT 13.800 127.100 14.600 127.200 ;
        RECT 15.900 127.100 16.200 127.800 ;
        RECT 20.700 127.700 21.100 127.800 ;
        RECT 22.200 127.700 22.600 129.900 ;
        RECT 20.700 127.400 22.600 127.700 ;
        RECT 18.700 127.100 19.100 127.200 ;
        RECT 12.600 126.800 19.300 127.100 ;
        RECT 15.300 126.700 15.700 126.800 ;
        RECT 10.200 125.800 12.200 126.100 ;
        RECT 14.500 126.200 14.900 126.300 ;
        RECT 15.800 126.200 16.200 126.300 ;
        RECT 14.500 125.900 17.000 126.200 ;
        RECT 16.600 125.800 17.000 125.900 ;
        RECT 10.200 125.400 10.600 125.800 ;
        RECT 9.100 124.600 9.900 124.900 ;
        RECT 7.000 121.500 7.400 123.500 ;
        RECT 9.100 121.100 9.500 124.600 ;
        RECT 11.800 121.100 12.200 125.800 ;
        RECT 13.400 125.500 16.200 125.600 ;
        RECT 13.400 125.400 16.300 125.500 ;
        RECT 13.400 125.300 18.300 125.400 ;
        RECT 13.400 121.100 13.800 125.300 ;
        RECT 15.900 125.100 18.300 125.300 ;
        RECT 15.000 124.500 17.700 124.800 ;
        RECT 15.000 124.400 15.400 124.500 ;
        RECT 17.300 124.400 17.700 124.500 ;
        RECT 18.000 124.500 18.300 125.100 ;
        RECT 19.000 125.200 19.300 126.800 ;
        RECT 19.800 126.400 20.200 126.500 ;
        RECT 19.800 126.100 21.700 126.400 ;
        RECT 21.300 126.000 21.700 126.100 ;
        RECT 20.500 125.700 20.900 125.800 ;
        RECT 22.200 125.700 22.600 127.400 ;
        RECT 24.800 127.100 25.200 129.900 ;
        RECT 26.200 127.500 26.600 129.900 ;
        RECT 28.400 129.200 28.800 129.900 ;
        RECT 27.800 128.900 28.800 129.200 ;
        RECT 30.600 128.900 31.000 129.900 ;
        RECT 32.700 129.200 33.300 129.900 ;
        RECT 32.600 128.900 33.300 129.200 ;
        RECT 27.800 128.500 28.200 128.900 ;
        RECT 30.600 128.600 30.900 128.900 ;
        RECT 28.600 128.200 29.000 128.600 ;
        RECT 29.500 128.300 30.900 128.600 ;
        RECT 32.600 128.500 33.000 128.900 ;
        RECT 29.500 128.200 29.900 128.300 ;
        RECT 26.600 127.100 27.400 127.200 ;
        RECT 28.700 127.100 29.000 128.200 ;
        RECT 33.500 127.700 33.900 127.800 ;
        RECT 35.000 127.700 35.400 129.900 ;
        RECT 33.500 127.400 35.400 127.700 ;
        RECT 31.500 127.100 31.900 127.200 ;
        RECT 24.800 126.900 25.700 127.100 ;
        RECT 24.900 126.800 25.700 126.900 ;
        RECT 26.600 126.800 32.100 127.100 ;
        RECT 23.800 125.800 24.600 126.200 ;
        RECT 20.500 125.400 22.600 125.700 ;
        RECT 19.000 124.900 20.200 125.200 ;
        RECT 18.700 124.500 19.100 124.600 ;
        RECT 18.000 124.200 19.100 124.500 ;
        RECT 19.900 124.400 20.200 124.900 ;
        RECT 20.600 124.800 21.000 125.400 ;
        RECT 19.900 124.000 20.600 124.400 ;
        RECT 16.700 123.700 17.100 123.800 ;
        RECT 18.100 123.700 18.500 123.800 ;
        RECT 15.000 123.100 15.400 123.500 ;
        RECT 16.700 123.400 18.500 123.700 ;
        RECT 17.800 123.100 18.100 123.400 ;
        RECT 19.800 123.100 20.200 123.500 ;
        RECT 15.000 122.800 16.000 123.100 ;
        RECT 15.600 121.100 16.000 122.800 ;
        RECT 17.800 121.100 18.200 123.100 ;
        RECT 19.900 121.100 20.500 123.100 ;
        RECT 22.200 121.100 22.600 125.400 ;
        RECT 23.000 124.800 23.400 125.600 ;
        RECT 25.400 125.200 25.700 126.800 ;
        RECT 28.100 126.700 28.500 126.800 ;
        RECT 27.300 126.200 27.700 126.300 ;
        RECT 27.300 125.900 29.800 126.200 ;
        RECT 29.400 125.800 29.800 125.900 ;
        RECT 26.200 125.500 29.000 125.600 ;
        RECT 26.200 125.400 29.100 125.500 ;
        RECT 26.200 125.300 31.100 125.400 ;
        RECT 25.400 124.800 25.800 125.200 ;
        RECT 24.600 123.800 25.000 124.600 ;
        RECT 25.400 123.500 25.700 124.800 ;
        RECT 23.900 123.200 25.700 123.500 ;
        RECT 23.900 123.100 24.200 123.200 ;
        RECT 23.800 121.100 24.200 123.100 ;
        RECT 25.400 123.100 25.700 123.200 ;
        RECT 25.400 121.100 25.800 123.100 ;
        RECT 26.200 121.100 26.600 125.300 ;
        RECT 28.700 125.100 31.100 125.300 ;
        RECT 27.800 124.500 30.500 124.800 ;
        RECT 27.800 124.400 28.200 124.500 ;
        RECT 30.100 124.400 30.500 124.500 ;
        RECT 30.800 124.500 31.100 125.100 ;
        RECT 31.800 125.200 32.100 126.800 ;
        RECT 32.600 126.400 33.000 126.500 ;
        RECT 32.600 126.100 34.500 126.400 ;
        RECT 34.100 126.000 34.500 126.100 ;
        RECT 33.300 125.700 33.700 125.800 ;
        RECT 35.000 125.700 35.400 127.400 ;
        RECT 37.400 128.500 37.800 129.500 ;
        RECT 37.400 127.400 37.700 128.500 ;
        RECT 39.500 128.200 39.900 129.500 ;
        RECT 39.000 128.000 39.900 128.200 ;
        RECT 39.000 127.800 40.300 128.000 ;
        RECT 39.500 127.700 40.300 127.800 ;
        RECT 39.900 127.500 40.300 127.700 ;
        RECT 37.400 127.100 39.500 127.400 ;
        RECT 39.000 126.900 39.500 127.100 ;
        RECT 40.000 127.200 40.300 127.500 ;
        RECT 37.400 125.800 37.800 126.600 ;
        RECT 38.200 125.800 38.600 126.600 ;
        RECT 39.000 126.500 39.700 126.900 ;
        RECT 40.000 126.800 41.000 127.200 ;
        RECT 33.300 125.400 35.400 125.700 ;
        RECT 39.000 125.500 39.300 126.500 ;
        RECT 31.800 124.900 33.000 125.200 ;
        RECT 31.500 124.500 31.900 124.600 ;
        RECT 30.800 124.200 31.900 124.500 ;
        RECT 32.700 124.400 33.000 124.900 ;
        RECT 32.700 124.000 33.400 124.400 ;
        RECT 29.500 123.700 29.900 123.800 ;
        RECT 30.900 123.700 31.300 123.800 ;
        RECT 27.800 123.100 28.200 123.500 ;
        RECT 29.500 123.400 31.300 123.700 ;
        RECT 30.600 123.100 30.900 123.400 ;
        RECT 32.600 123.100 33.000 123.500 ;
        RECT 27.800 122.800 28.800 123.100 ;
        RECT 28.400 121.100 28.800 122.800 ;
        RECT 30.600 121.100 31.000 123.100 ;
        RECT 32.700 121.100 33.300 123.100 ;
        RECT 35.000 121.100 35.400 125.400 ;
        RECT 37.400 125.200 39.300 125.500 ;
        RECT 37.400 123.500 37.700 125.200 ;
        RECT 40.000 124.900 40.300 126.800 ;
        RECT 40.600 126.100 41.000 126.200 ;
        RECT 42.200 126.100 42.600 129.900 ;
        RECT 43.000 127.800 43.400 128.600 ;
        RECT 43.800 128.500 44.200 129.500 ;
        RECT 43.800 127.400 44.100 128.500 ;
        RECT 45.900 128.200 46.300 129.500 ;
        RECT 45.400 128.000 46.300 128.200 ;
        RECT 45.400 127.800 46.700 128.000 ;
        RECT 45.900 127.700 46.700 127.800 ;
        RECT 46.300 127.500 46.700 127.700 ;
        RECT 43.800 127.100 45.900 127.400 ;
        RECT 45.400 126.900 45.900 127.100 ;
        RECT 46.400 127.200 46.700 127.500 ;
        RECT 40.600 125.800 42.600 126.100 ;
        RECT 43.800 125.800 44.200 126.600 ;
        RECT 44.600 125.800 45.000 126.600 ;
        RECT 45.400 126.500 46.100 126.900 ;
        RECT 46.400 126.800 47.400 127.200 ;
        RECT 40.600 125.400 41.000 125.800 ;
        RECT 39.500 124.600 40.300 124.900 ;
        RECT 37.400 121.500 37.800 123.500 ;
        RECT 39.500 121.100 39.900 124.600 ;
        RECT 42.200 121.100 42.600 125.800 ;
        RECT 45.400 125.500 45.700 126.500 ;
        RECT 43.800 125.200 45.700 125.500 ;
        RECT 43.800 123.500 44.100 125.200 ;
        RECT 46.400 124.900 46.700 126.800 ;
        RECT 47.000 126.100 47.400 126.200 ;
        RECT 48.600 126.100 49.000 129.900 ;
        RECT 49.400 127.800 49.800 128.600 ;
        RECT 50.200 127.500 50.600 129.900 ;
        RECT 52.400 129.200 52.800 129.900 ;
        RECT 51.800 128.900 52.800 129.200 ;
        RECT 54.600 128.900 55.000 129.900 ;
        RECT 56.700 129.200 57.300 129.900 ;
        RECT 56.600 128.900 57.300 129.200 ;
        RECT 51.800 128.500 52.200 128.900 ;
        RECT 54.600 128.600 54.900 128.900 ;
        RECT 52.600 127.800 53.000 128.600 ;
        RECT 53.500 128.300 54.900 128.600 ;
        RECT 56.600 128.500 57.000 128.900 ;
        RECT 53.500 128.200 53.900 128.300 ;
        RECT 50.600 127.100 51.400 127.200 ;
        RECT 52.700 127.100 53.000 127.800 ;
        RECT 57.500 127.700 57.900 127.800 ;
        RECT 59.000 127.700 59.400 129.900 ;
        RECT 57.500 127.400 59.400 127.700 ;
        RECT 55.500 127.100 55.900 127.200 ;
        RECT 50.600 126.800 56.100 127.100 ;
        RECT 52.100 126.700 52.500 126.800 ;
        RECT 47.000 125.800 49.000 126.100 ;
        RECT 51.300 126.200 51.700 126.300 ;
        RECT 51.300 125.900 53.800 126.200 ;
        RECT 53.400 125.800 53.800 125.900 ;
        RECT 47.000 125.400 47.400 125.800 ;
        RECT 45.900 124.600 46.700 124.900 ;
        RECT 43.800 121.500 44.200 123.500 ;
        RECT 45.900 121.100 46.300 124.600 ;
        RECT 48.600 121.100 49.000 125.800 ;
        RECT 50.200 125.500 53.000 125.600 ;
        RECT 50.200 125.400 53.100 125.500 ;
        RECT 50.200 125.300 55.100 125.400 ;
        RECT 50.200 121.100 50.600 125.300 ;
        RECT 52.700 125.100 55.100 125.300 ;
        RECT 51.800 124.500 54.500 124.800 ;
        RECT 51.800 124.400 52.200 124.500 ;
        RECT 54.100 124.400 54.500 124.500 ;
        RECT 54.800 124.500 55.100 125.100 ;
        RECT 55.800 125.200 56.100 126.800 ;
        RECT 56.600 126.400 57.000 126.500 ;
        RECT 56.600 126.100 58.500 126.400 ;
        RECT 58.100 126.000 58.500 126.100 ;
        RECT 57.300 125.700 57.700 125.800 ;
        RECT 59.000 125.700 59.400 127.400 ;
        RECT 60.400 128.200 60.800 129.900 ;
        RECT 60.400 127.800 61.000 128.200 ;
        RECT 60.400 127.100 60.800 127.800 ;
        RECT 57.300 125.400 59.400 125.700 ;
        RECT 55.800 124.900 57.000 125.200 ;
        RECT 55.500 124.500 55.900 124.600 ;
        RECT 54.800 124.200 55.900 124.500 ;
        RECT 56.700 124.400 57.000 124.900 ;
        RECT 56.700 124.000 57.400 124.400 ;
        RECT 53.500 123.700 53.900 123.800 ;
        RECT 54.900 123.700 55.300 123.800 ;
        RECT 51.800 123.100 52.200 123.500 ;
        RECT 53.500 123.400 55.300 123.700 ;
        RECT 54.600 123.100 54.900 123.400 ;
        RECT 56.600 123.100 57.000 123.500 ;
        RECT 51.800 122.800 52.800 123.100 ;
        RECT 52.400 121.100 52.800 122.800 ;
        RECT 54.600 121.100 55.000 123.100 ;
        RECT 56.700 121.100 57.300 123.100 ;
        RECT 59.000 121.100 59.400 125.400 ;
        RECT 59.900 126.900 60.800 127.100 ;
        RECT 64.800 127.100 65.200 129.900 ;
        RECT 66.800 127.100 67.200 129.900 ;
        RECT 64.800 126.900 65.700 127.100 ;
        RECT 59.900 126.800 60.700 126.900 ;
        RECT 64.900 126.800 65.700 126.900 ;
        RECT 59.900 125.200 60.200 126.800 ;
        RECT 65.400 126.200 65.700 126.800 ;
        RECT 66.300 126.900 67.200 127.100 ;
        RECT 71.200 127.100 71.600 129.900 ;
        RECT 74.400 127.100 74.800 129.900 ;
        RECT 77.400 129.200 77.800 129.900 ;
        RECT 79.000 129.200 79.400 129.900 ;
        RECT 77.400 128.900 77.900 129.200 ;
        RECT 77.600 128.800 77.900 128.900 ;
        RECT 79.000 128.800 80.200 129.200 ;
        RECT 77.600 128.500 79.600 128.800 ;
        RECT 75.800 128.100 76.200 128.200 ;
        RECT 76.600 128.100 77.500 128.200 ;
        RECT 75.800 127.800 77.500 128.100 ;
        RECT 76.600 127.100 77.000 127.200 ;
        RECT 77.400 127.100 78.200 127.200 ;
        RECT 71.200 126.900 72.100 127.100 ;
        RECT 74.400 126.900 75.300 127.100 ;
        RECT 66.300 126.800 67.100 126.900 ;
        RECT 71.300 126.800 72.100 126.900 ;
        RECT 74.500 126.800 75.300 126.900 ;
        RECT 76.600 126.800 78.200 127.100 ;
        RECT 61.000 125.800 61.800 126.200 ;
        RECT 63.800 125.800 64.600 126.200 ;
        RECT 65.400 125.800 65.800 126.200 ;
        RECT 59.800 124.800 60.200 125.200 ;
        RECT 62.200 124.800 62.600 125.600 ;
        RECT 63.000 124.800 63.400 125.600 ;
        RECT 65.400 125.200 65.700 125.800 ;
        RECT 66.300 125.200 66.600 126.800 ;
        RECT 67.400 125.800 68.200 126.200 ;
        RECT 70.200 125.800 71.000 126.200 ;
        RECT 65.400 124.800 65.800 125.200 ;
        RECT 66.200 124.800 66.600 125.200 ;
        RECT 68.600 124.800 69.000 125.600 ;
        RECT 69.400 124.800 69.800 125.600 ;
        RECT 71.800 125.200 72.100 126.800 ;
        RECT 73.400 125.800 74.200 126.200 ;
        RECT 71.800 124.800 72.200 125.200 ;
        RECT 72.600 124.800 73.000 125.600 ;
        RECT 75.000 125.200 75.300 126.800 ;
        RECT 78.200 125.800 79.000 126.200 ;
        RECT 79.300 125.200 79.600 128.500 ;
        RECT 82.200 127.500 82.600 129.900 ;
        RECT 84.400 129.200 84.800 129.900 ;
        RECT 83.800 128.900 84.800 129.200 ;
        RECT 86.600 128.900 87.000 129.900 ;
        RECT 88.700 129.200 89.300 129.900 ;
        RECT 88.600 128.900 89.300 129.200 ;
        RECT 83.800 128.500 84.200 128.900 ;
        RECT 86.600 128.600 86.900 128.900 ;
        RECT 84.600 128.200 85.000 128.600 ;
        RECT 85.500 128.300 86.900 128.600 ;
        RECT 88.600 128.500 89.000 128.900 ;
        RECT 85.500 128.200 85.900 128.300 ;
        RECT 82.600 127.100 83.400 127.200 ;
        RECT 84.700 127.100 85.000 128.200 ;
        RECT 91.000 128.100 91.400 129.900 ;
        RECT 93.400 128.100 93.800 128.600 ;
        RECT 91.000 127.800 93.800 128.100 ;
        RECT 89.500 127.700 89.900 127.800 ;
        RECT 91.000 127.700 91.400 127.800 ;
        RECT 89.500 127.400 91.400 127.700 ;
        RECT 85.400 127.100 85.800 127.200 ;
        RECT 87.500 127.100 87.900 127.200 ;
        RECT 82.600 126.800 88.100 127.100 ;
        RECT 84.100 126.700 84.500 126.800 ;
        RECT 83.300 126.200 83.700 126.300 ;
        RECT 83.300 126.100 85.800 126.200 ;
        RECT 86.200 126.100 86.600 126.200 ;
        RECT 83.300 125.900 86.600 126.100 ;
        RECT 85.400 125.800 86.600 125.900 ;
        RECT 82.200 125.500 85.000 125.600 ;
        RECT 82.200 125.400 85.100 125.500 ;
        RECT 82.200 125.300 87.100 125.400 ;
        RECT 75.000 124.800 75.400 125.200 ;
        RECT 79.300 124.900 81.000 125.200 ;
        RECT 80.600 124.800 81.000 124.900 ;
        RECT 59.900 123.500 60.200 124.800 ;
        RECT 60.600 123.800 61.000 124.600 ;
        RECT 64.600 123.800 65.000 124.600 ;
        RECT 65.400 123.500 65.700 124.800 ;
        RECT 59.900 123.200 61.700 123.500 ;
        RECT 59.900 123.100 60.200 123.200 ;
        RECT 59.800 121.100 60.200 123.100 ;
        RECT 61.400 123.100 61.700 123.200 ;
        RECT 63.900 123.200 65.700 123.500 ;
        RECT 63.900 123.100 64.200 123.200 ;
        RECT 61.400 121.100 61.800 123.100 ;
        RECT 63.800 121.100 64.200 123.100 ;
        RECT 65.400 123.100 65.700 123.200 ;
        RECT 66.300 123.500 66.600 124.800 ;
        RECT 67.000 123.800 67.400 124.600 ;
        RECT 69.400 124.100 69.700 124.800 ;
        RECT 67.800 123.800 69.700 124.100 ;
        RECT 71.000 123.800 71.400 124.600 ;
        RECT 67.800 123.500 68.100 123.800 ;
        RECT 71.800 123.500 72.100 124.800 ;
        RECT 74.200 123.800 74.600 124.600 ;
        RECT 75.000 123.500 75.300 124.800 ;
        RECT 75.900 124.400 77.700 124.700 ;
        RECT 75.900 124.100 76.200 124.400 ;
        RECT 66.300 123.200 68.100 123.500 ;
        RECT 66.300 123.100 66.600 123.200 ;
        RECT 65.400 121.100 65.800 123.100 ;
        RECT 66.200 121.100 66.600 123.100 ;
        RECT 67.800 123.100 68.100 123.200 ;
        RECT 70.300 123.200 72.100 123.500 ;
        RECT 70.300 123.100 70.600 123.200 ;
        RECT 67.800 121.100 68.200 123.100 ;
        RECT 70.200 121.100 70.600 123.100 ;
        RECT 71.800 123.100 72.100 123.200 ;
        RECT 73.500 123.200 75.300 123.500 ;
        RECT 73.500 123.100 73.800 123.200 ;
        RECT 71.800 121.100 72.200 123.100 ;
        RECT 73.400 121.100 73.800 123.100 ;
        RECT 75.000 123.100 75.300 123.200 ;
        RECT 75.000 121.100 75.400 123.100 ;
        RECT 75.800 121.100 76.200 124.100 ;
        RECT 77.400 124.100 77.700 124.400 ;
        RECT 78.300 124.500 80.100 124.600 ;
        RECT 80.600 124.500 80.900 124.800 ;
        RECT 78.300 124.300 80.200 124.500 ;
        RECT 78.300 124.100 78.600 124.300 ;
        RECT 77.400 121.400 77.800 124.100 ;
        RECT 78.200 121.700 78.600 124.100 ;
        RECT 79.000 121.400 79.400 124.000 ;
        RECT 79.800 121.500 80.200 124.300 ;
        RECT 80.600 121.700 81.000 124.500 ;
        RECT 77.400 121.100 79.400 121.400 ;
        RECT 79.900 121.400 80.200 121.500 ;
        RECT 81.400 121.500 81.800 124.500 ;
        RECT 81.400 121.400 81.700 121.500 ;
        RECT 79.900 121.100 81.700 121.400 ;
        RECT 82.200 121.100 82.600 125.300 ;
        RECT 84.700 125.100 87.100 125.300 ;
        RECT 83.800 124.500 86.500 124.800 ;
        RECT 83.800 124.400 84.200 124.500 ;
        RECT 86.100 124.400 86.500 124.500 ;
        RECT 86.800 124.500 87.100 125.100 ;
        RECT 87.800 125.200 88.100 126.800 ;
        RECT 88.600 126.400 89.000 126.500 ;
        RECT 88.600 126.100 90.500 126.400 ;
        RECT 90.100 126.000 90.500 126.100 ;
        RECT 89.300 125.700 89.700 125.800 ;
        RECT 91.000 125.700 91.400 127.400 ;
        RECT 89.300 125.400 91.400 125.700 ;
        RECT 87.800 124.900 89.000 125.200 ;
        RECT 87.500 124.500 87.900 124.600 ;
        RECT 86.800 124.200 87.900 124.500 ;
        RECT 88.700 124.400 89.000 124.900 ;
        RECT 88.700 124.000 89.400 124.400 ;
        RECT 91.000 124.100 91.400 125.400 ;
        RECT 94.200 126.100 94.600 129.900 ;
        RECT 96.900 128.000 97.300 129.500 ;
        RECT 99.000 128.500 99.400 129.500 ;
        RECT 96.500 127.700 97.300 128.000 ;
        RECT 96.500 127.500 96.900 127.700 ;
        RECT 96.500 127.200 96.800 127.500 ;
        RECT 99.100 127.400 99.400 128.500 ;
        RECT 100.100 128.200 100.500 129.900 ;
        RECT 100.100 127.900 101.000 128.200 ;
        RECT 95.000 127.100 95.400 127.200 ;
        RECT 95.800 127.100 96.800 127.200 ;
        RECT 95.000 126.800 96.800 127.100 ;
        RECT 97.300 127.100 99.400 127.400 ;
        RECT 97.300 126.900 97.800 127.100 ;
        RECT 95.800 126.100 96.200 126.200 ;
        RECT 94.200 125.800 96.200 126.100 ;
        RECT 93.400 124.100 93.800 124.200 ;
        RECT 91.000 123.800 93.800 124.100 ;
        RECT 85.500 123.700 85.900 123.800 ;
        RECT 86.900 123.700 87.300 123.800 ;
        RECT 83.800 123.100 84.200 123.500 ;
        RECT 85.500 123.400 87.300 123.700 ;
        RECT 86.600 123.100 86.900 123.400 ;
        RECT 88.600 123.100 89.000 123.500 ;
        RECT 83.800 122.800 84.800 123.100 ;
        RECT 84.400 121.100 84.800 122.800 ;
        RECT 86.600 121.100 87.000 123.100 ;
        RECT 88.700 121.100 89.300 123.100 ;
        RECT 91.000 121.100 91.400 123.800 ;
        RECT 94.200 121.100 94.600 125.800 ;
        RECT 95.800 125.400 96.200 125.800 ;
        RECT 96.500 124.900 96.800 126.800 ;
        RECT 97.100 126.500 97.800 126.900 ;
        RECT 99.800 126.800 100.200 127.200 ;
        RECT 97.500 125.500 97.800 126.500 ;
        RECT 98.200 125.800 98.600 126.600 ;
        RECT 99.000 125.800 99.400 126.600 ;
        RECT 99.800 126.100 100.100 126.800 ;
        RECT 100.600 126.100 101.000 127.900 ;
        RECT 103.800 127.900 104.200 129.900 ;
        RECT 106.200 128.900 106.600 129.900 ;
        RECT 104.500 128.200 104.900 128.600 ;
        RECT 104.600 128.100 105.000 128.200 ;
        RECT 106.200 128.100 106.500 128.900 ;
        RECT 101.400 126.800 101.800 127.600 ;
        RECT 103.000 126.400 103.400 127.200 ;
        RECT 99.800 125.800 101.000 126.100 ;
        RECT 102.200 126.100 102.600 126.200 ;
        RECT 103.800 126.100 104.100 127.900 ;
        RECT 104.600 127.800 106.500 128.100 ;
        RECT 107.000 127.800 107.400 128.600 ;
        RECT 106.200 127.200 106.500 127.800 ;
        RECT 107.800 127.700 108.200 129.900 ;
        RECT 109.900 129.200 110.500 129.900 ;
        RECT 109.900 128.900 110.600 129.200 ;
        RECT 112.200 128.900 112.600 129.900 ;
        RECT 114.400 129.200 114.800 129.900 ;
        RECT 114.400 128.900 115.400 129.200 ;
        RECT 110.200 128.500 110.600 128.900 ;
        RECT 112.300 128.600 112.600 128.900 ;
        RECT 112.300 128.300 113.700 128.600 ;
        RECT 113.300 128.200 113.700 128.300 ;
        RECT 114.200 128.200 114.600 128.600 ;
        RECT 115.000 128.500 115.400 128.900 ;
        RECT 109.300 127.700 109.700 127.800 ;
        RECT 107.800 127.400 109.700 127.700 ;
        RECT 106.200 126.800 106.600 127.200 ;
        RECT 104.600 126.100 105.000 126.200 ;
        RECT 102.200 125.800 103.000 126.100 ;
        RECT 103.800 125.800 105.000 126.100 ;
        RECT 97.500 125.200 99.400 125.500 ;
        RECT 96.500 124.600 97.300 124.900 ;
        RECT 96.900 121.100 97.300 124.600 ;
        RECT 99.100 123.500 99.400 125.200 ;
        RECT 99.800 124.400 100.200 125.200 ;
        RECT 99.000 121.500 99.400 123.500 ;
        RECT 100.600 121.100 101.000 125.800 ;
        RECT 102.600 125.600 103.000 125.800 ;
        RECT 104.600 125.100 104.900 125.800 ;
        RECT 105.400 125.400 105.800 126.200 ;
        RECT 106.200 125.100 106.500 126.800 ;
        RECT 107.800 125.700 108.200 127.400 ;
        RECT 111.300 127.100 111.700 127.200 ;
        RECT 114.200 127.100 114.500 128.200 ;
        RECT 116.600 127.500 117.000 129.900 ;
        RECT 117.400 127.700 117.800 129.900 ;
        RECT 119.500 129.200 120.100 129.900 ;
        RECT 119.500 128.900 120.200 129.200 ;
        RECT 121.800 128.900 122.200 129.900 ;
        RECT 124.000 129.200 124.400 129.900 ;
        RECT 124.000 128.900 125.000 129.200 ;
        RECT 119.800 128.500 120.200 128.900 ;
        RECT 121.900 128.600 122.200 128.900 ;
        RECT 121.900 128.300 123.300 128.600 ;
        RECT 122.900 128.200 123.300 128.300 ;
        RECT 120.600 127.800 121.000 128.200 ;
        RECT 123.800 127.800 124.200 128.600 ;
        RECT 124.600 128.500 125.000 128.900 ;
        RECT 118.900 127.700 119.300 127.800 ;
        RECT 117.400 127.400 119.300 127.700 ;
        RECT 115.800 127.100 116.600 127.200 ;
        RECT 111.100 126.800 116.600 127.100 ;
        RECT 110.200 126.400 110.600 126.500 ;
        RECT 108.700 126.100 110.600 126.400 ;
        RECT 108.700 126.000 109.100 126.100 ;
        RECT 109.500 125.700 109.900 125.800 ;
        RECT 107.800 125.400 109.900 125.700 ;
        RECT 102.200 124.800 104.200 125.100 ;
        RECT 102.200 121.100 102.600 124.800 ;
        RECT 103.800 121.100 104.200 124.800 ;
        RECT 104.600 121.100 105.000 125.100 ;
        RECT 105.700 124.700 106.600 125.100 ;
        RECT 105.700 121.100 106.100 124.700 ;
        RECT 107.800 121.100 108.200 125.400 ;
        RECT 111.100 125.200 111.400 126.800 ;
        RECT 114.700 126.700 115.100 126.800 ;
        RECT 115.500 126.200 115.900 126.300 ;
        RECT 113.400 125.900 115.900 126.200 ;
        RECT 113.400 125.800 113.800 125.900 ;
        RECT 117.400 125.700 117.800 127.400 ;
        RECT 120.600 127.200 120.900 127.800 ;
        RECT 120.600 127.100 121.300 127.200 ;
        RECT 123.800 127.100 124.100 127.800 ;
        RECT 126.200 127.500 126.600 129.900 ;
        RECT 127.000 127.800 127.400 128.600 ;
        RECT 125.400 127.100 126.200 127.200 ;
        RECT 120.600 126.800 126.200 127.100 ;
        RECT 127.000 127.100 127.400 127.200 ;
        RECT 127.800 127.100 128.200 129.900 ;
        RECT 133.400 129.600 135.400 129.900 ;
        RECT 128.600 128.500 129.000 129.500 ;
        RECT 128.600 127.400 128.900 128.500 ;
        RECT 130.700 128.200 131.100 129.500 ;
        RECT 130.200 128.000 131.100 128.200 ;
        RECT 130.200 127.800 131.500 128.000 ;
        RECT 133.400 127.900 133.800 129.600 ;
        RECT 134.200 127.900 134.600 129.300 ;
        RECT 135.000 128.000 135.400 129.600 ;
        RECT 136.600 128.000 137.000 129.900 ;
        RECT 135.000 127.900 137.000 128.000 ;
        RECT 130.700 127.700 131.500 127.800 ;
        RECT 131.100 127.500 131.500 127.700 ;
        RECT 128.600 127.100 130.700 127.400 ;
        RECT 127.000 126.800 128.200 127.100 ;
        RECT 119.800 126.400 120.200 126.500 ;
        RECT 118.300 126.100 120.200 126.400 ;
        RECT 118.300 126.000 118.700 126.100 ;
        RECT 119.100 125.700 119.500 125.800 ;
        RECT 114.200 125.500 117.000 125.600 ;
        RECT 114.100 125.400 117.000 125.500 ;
        RECT 110.200 124.900 111.400 125.200 ;
        RECT 112.100 125.300 117.000 125.400 ;
        RECT 112.100 125.100 114.500 125.300 ;
        RECT 110.200 124.400 110.500 124.900 ;
        RECT 109.800 124.000 110.500 124.400 ;
        RECT 111.300 124.500 111.700 124.600 ;
        RECT 112.100 124.500 112.400 125.100 ;
        RECT 111.300 124.200 112.400 124.500 ;
        RECT 112.700 124.500 115.400 124.800 ;
        RECT 112.700 124.400 113.100 124.500 ;
        RECT 115.000 124.400 115.400 124.500 ;
        RECT 111.900 123.700 112.300 123.800 ;
        RECT 113.300 123.700 113.700 123.800 ;
        RECT 110.200 123.100 110.600 123.500 ;
        RECT 111.900 123.400 113.700 123.700 ;
        RECT 112.300 123.100 112.600 123.400 ;
        RECT 115.000 123.100 115.400 123.500 ;
        RECT 109.900 121.100 110.500 123.100 ;
        RECT 112.200 121.100 112.600 123.100 ;
        RECT 114.400 122.800 115.400 123.100 ;
        RECT 114.400 121.100 114.800 122.800 ;
        RECT 116.600 121.100 117.000 125.300 ;
        RECT 117.400 125.400 119.500 125.700 ;
        RECT 117.400 121.100 117.800 125.400 ;
        RECT 120.700 125.200 121.000 126.800 ;
        RECT 124.300 126.700 124.700 126.800 ;
        RECT 123.800 126.200 124.200 126.300 ;
        RECT 125.100 126.200 125.500 126.300 ;
        RECT 123.000 125.900 125.500 126.200 ;
        RECT 123.000 125.800 123.400 125.900 ;
        RECT 123.800 125.500 126.600 125.600 ;
        RECT 123.700 125.400 126.600 125.500 ;
        RECT 119.800 124.900 121.000 125.200 ;
        RECT 121.700 125.300 126.600 125.400 ;
        RECT 121.700 125.100 124.100 125.300 ;
        RECT 119.800 124.400 120.100 124.900 ;
        RECT 119.400 124.000 120.100 124.400 ;
        RECT 120.900 124.500 121.300 124.600 ;
        RECT 121.700 124.500 122.000 125.100 ;
        RECT 120.900 124.200 122.000 124.500 ;
        RECT 122.300 124.500 125.000 124.800 ;
        RECT 122.300 124.400 122.700 124.500 ;
        RECT 124.600 124.400 125.000 124.500 ;
        RECT 121.500 123.700 121.900 123.800 ;
        RECT 122.900 123.700 123.300 123.800 ;
        RECT 119.800 123.100 120.200 123.500 ;
        RECT 121.500 123.400 123.300 123.700 ;
        RECT 121.900 123.100 122.200 123.400 ;
        RECT 124.600 123.100 125.000 123.500 ;
        RECT 119.500 121.100 120.100 123.100 ;
        RECT 121.800 121.100 122.200 123.100 ;
        RECT 124.000 122.800 125.000 123.100 ;
        RECT 124.000 121.100 124.400 122.800 ;
        RECT 126.200 121.100 126.600 125.300 ;
        RECT 127.800 121.100 128.200 126.800 ;
        RECT 130.200 126.900 130.700 127.100 ;
        RECT 131.200 127.200 131.500 127.500 ;
        RECT 134.200 127.200 134.500 127.900 ;
        RECT 135.100 127.700 136.900 127.900 ;
        RECT 136.200 127.200 136.600 127.400 ;
        RECT 128.600 125.800 129.000 126.600 ;
        RECT 129.400 125.800 129.800 126.600 ;
        RECT 130.200 126.500 130.900 126.900 ;
        RECT 131.200 126.800 132.200 127.200 ;
        RECT 130.200 125.500 130.500 126.500 ;
        RECT 128.600 125.200 130.500 125.500 ;
        RECT 128.600 123.500 128.900 125.200 ;
        RECT 131.200 124.900 131.500 126.800 ;
        RECT 133.400 126.400 133.800 127.200 ;
        RECT 134.200 126.900 135.400 127.200 ;
        RECT 136.200 127.100 137.000 127.200 ;
        RECT 137.400 127.100 137.800 129.900 ;
        RECT 138.200 128.100 138.600 128.600 ;
        RECT 139.000 128.100 139.400 128.200 ;
        RECT 138.200 127.800 139.400 128.100 ;
        RECT 142.200 127.900 142.600 129.900 ;
        RECT 146.200 128.900 146.600 129.900 ;
        RECT 147.800 129.200 148.200 129.900 ;
        RECT 146.000 128.800 146.600 128.900 ;
        RECT 147.700 128.800 148.200 129.200 ;
        RECT 142.900 128.200 143.300 128.600 ;
        RECT 146.000 128.500 148.000 128.800 ;
        RECT 136.200 126.900 137.800 127.100 ;
        RECT 135.000 126.800 135.400 126.900 ;
        RECT 136.600 126.800 137.800 126.900 ;
        RECT 140.600 127.100 141.000 127.200 ;
        RECT 141.400 127.100 141.800 127.200 ;
        RECT 140.600 126.800 141.800 127.100 ;
        RECT 131.800 125.400 132.200 126.200 ;
        RECT 134.200 125.800 134.600 126.600 ;
        RECT 135.100 125.100 135.400 126.800 ;
        RECT 135.800 125.800 136.200 126.600 ;
        RECT 130.700 124.600 131.500 124.900 ;
        RECT 128.600 121.500 129.000 123.500 ;
        RECT 130.700 121.100 131.100 124.600 ;
        RECT 134.700 121.100 135.700 125.100 ;
        RECT 137.400 121.100 137.800 126.800 ;
        RECT 141.400 126.400 141.800 126.800 ;
        RECT 140.600 126.100 141.000 126.200 ;
        RECT 142.200 126.100 142.500 127.900 ;
        RECT 143.000 127.800 143.400 128.200 ;
        RECT 143.000 126.100 143.400 126.200 ;
        RECT 140.600 125.800 141.400 126.100 ;
        RECT 142.200 125.800 143.400 126.100 ;
        RECT 141.000 125.600 141.400 125.800 ;
        RECT 143.000 125.100 143.300 125.800 ;
        RECT 146.000 125.200 146.300 128.500 ;
        RECT 148.100 128.100 149.000 128.200 ;
        RECT 149.400 128.100 149.800 128.200 ;
        RECT 148.100 127.800 149.800 128.100 ;
        RECT 150.200 127.700 150.600 129.900 ;
        RECT 152.300 129.200 152.900 129.900 ;
        RECT 152.300 128.900 153.000 129.200 ;
        RECT 154.600 128.900 155.000 129.900 ;
        RECT 156.800 129.200 157.200 129.900 ;
        RECT 156.800 128.900 157.800 129.200 ;
        RECT 152.600 128.500 153.000 128.900 ;
        RECT 154.700 128.600 155.000 128.900 ;
        RECT 154.700 128.300 156.100 128.600 ;
        RECT 155.700 128.200 156.100 128.300 ;
        RECT 156.600 128.200 157.000 128.600 ;
        RECT 157.400 128.500 157.800 128.900 ;
        RECT 151.700 127.700 152.100 127.800 ;
        RECT 150.200 127.400 152.100 127.700 ;
        RECT 147.400 127.100 148.200 127.200 ;
        RECT 148.600 127.100 149.000 127.200 ;
        RECT 147.400 126.800 149.000 127.100 ;
        RECT 146.600 125.800 147.400 126.200 ;
        RECT 140.600 124.800 142.600 125.100 ;
        RECT 140.600 121.100 141.000 124.800 ;
        RECT 142.200 121.100 142.600 124.800 ;
        RECT 143.000 121.100 143.400 125.100 ;
        RECT 144.600 124.900 146.300 125.200 ;
        RECT 150.200 125.700 150.600 127.400 ;
        RECT 153.700 127.100 154.100 127.200 ;
        RECT 155.800 127.100 156.200 127.200 ;
        RECT 156.600 127.100 156.900 128.200 ;
        RECT 159.000 127.500 159.400 129.900 ;
        RECT 159.800 129.600 161.800 129.900 ;
        RECT 159.800 127.900 160.200 129.600 ;
        RECT 160.600 127.900 161.000 129.300 ;
        RECT 161.400 128.000 161.800 129.600 ;
        RECT 163.000 128.000 163.400 129.900 ;
        RECT 161.400 127.900 163.400 128.000 ;
        RECT 163.800 128.500 164.200 129.500 ;
        RECT 160.600 127.200 160.900 127.900 ;
        RECT 161.500 127.700 163.300 127.900 ;
        RECT 163.800 127.400 164.100 128.500 ;
        RECT 165.900 128.000 166.300 129.500 ;
        RECT 169.400 128.900 169.800 129.900 ;
        RECT 165.900 127.700 166.700 128.000 ;
        RECT 166.300 127.500 166.700 127.700 ;
        RECT 162.600 127.200 163.000 127.400 ;
        RECT 158.200 127.100 159.000 127.200 ;
        RECT 153.500 126.800 159.000 127.100 ;
        RECT 152.600 126.400 153.000 126.500 ;
        RECT 151.100 126.100 153.000 126.400 ;
        RECT 153.500 126.200 153.800 126.800 ;
        RECT 157.100 126.700 157.500 126.800 ;
        RECT 159.800 126.400 160.200 127.200 ;
        RECT 160.600 126.900 161.800 127.200 ;
        RECT 162.600 126.900 163.400 127.200 ;
        RECT 163.800 127.100 165.900 127.400 ;
        RECT 161.400 126.800 161.800 126.900 ;
        RECT 163.000 126.800 163.400 126.900 ;
        RECT 165.400 126.900 165.900 127.100 ;
        RECT 166.400 127.200 166.700 127.500 ;
        RECT 169.400 127.200 169.700 128.900 ;
        RECT 170.200 127.800 170.600 128.600 ;
        RECT 171.000 127.500 171.400 129.900 ;
        RECT 173.200 129.200 173.600 129.900 ;
        RECT 172.600 128.900 173.600 129.200 ;
        RECT 175.400 128.900 175.800 129.900 ;
        RECT 177.500 129.200 178.100 129.900 ;
        RECT 177.400 128.900 178.100 129.200 ;
        RECT 172.600 128.500 173.000 128.900 ;
        RECT 175.400 128.600 175.700 128.900 ;
        RECT 173.400 128.200 173.800 128.600 ;
        RECT 174.300 128.300 175.700 128.600 ;
        RECT 177.400 128.500 177.800 128.900 ;
        RECT 174.300 128.200 174.700 128.300 ;
        RECT 157.900 126.200 158.300 126.300 ;
        RECT 151.100 126.000 151.500 126.100 ;
        RECT 153.400 125.800 153.800 126.200 ;
        RECT 155.000 126.100 155.400 126.200 ;
        RECT 155.800 126.100 158.300 126.200 ;
        RECT 155.000 125.900 158.300 126.100 ;
        RECT 155.000 125.800 156.200 125.900 ;
        RECT 160.600 125.800 161.000 126.600 ;
        RECT 151.900 125.700 152.300 125.800 ;
        RECT 150.200 125.400 152.300 125.700 ;
        RECT 144.600 124.800 145.000 124.900 ;
        RECT 144.700 124.500 145.000 124.800 ;
        RECT 145.500 124.500 147.300 124.600 ;
        RECT 143.800 121.500 144.200 124.500 ;
        RECT 144.600 121.700 145.000 124.500 ;
        RECT 145.400 124.300 147.300 124.500 ;
        RECT 143.900 121.400 144.200 121.500 ;
        RECT 145.400 121.500 145.800 124.300 ;
        RECT 147.000 124.100 147.300 124.300 ;
        RECT 147.900 124.400 149.700 124.700 ;
        RECT 147.900 124.100 148.200 124.400 ;
        RECT 145.400 121.400 145.700 121.500 ;
        RECT 143.900 121.100 145.700 121.400 ;
        RECT 146.200 121.400 146.600 124.000 ;
        RECT 147.000 121.700 147.400 124.100 ;
        RECT 147.800 121.400 148.200 124.100 ;
        RECT 146.200 121.100 148.200 121.400 ;
        RECT 149.400 124.100 149.700 124.400 ;
        RECT 149.400 121.100 149.800 124.100 ;
        RECT 150.200 121.100 150.600 125.400 ;
        RECT 153.500 125.200 153.800 125.800 ;
        RECT 156.600 125.500 159.400 125.600 ;
        RECT 156.500 125.400 159.400 125.500 ;
        RECT 152.600 124.900 153.800 125.200 ;
        RECT 154.500 125.300 159.400 125.400 ;
        RECT 154.500 125.100 156.900 125.300 ;
        RECT 152.600 124.400 152.900 124.900 ;
        RECT 152.200 124.000 152.900 124.400 ;
        RECT 153.700 124.500 154.100 124.600 ;
        RECT 154.500 124.500 154.800 125.100 ;
        RECT 153.700 124.200 154.800 124.500 ;
        RECT 155.100 124.500 157.800 124.800 ;
        RECT 155.100 124.400 155.500 124.500 ;
        RECT 157.400 124.400 157.800 124.500 ;
        RECT 154.300 123.700 154.700 123.800 ;
        RECT 155.700 123.700 156.100 123.800 ;
        RECT 152.600 123.100 153.000 123.500 ;
        RECT 154.300 123.400 156.100 123.700 ;
        RECT 154.700 123.100 155.000 123.400 ;
        RECT 157.400 123.100 157.800 123.500 ;
        RECT 152.300 121.100 152.900 123.100 ;
        RECT 154.600 121.100 155.000 123.100 ;
        RECT 156.800 122.800 157.800 123.100 ;
        RECT 156.800 121.100 157.200 122.800 ;
        RECT 159.000 121.100 159.400 125.300 ;
        RECT 161.500 125.100 161.800 126.800 ;
        RECT 162.200 125.800 162.600 126.600 ;
        RECT 163.000 126.100 163.400 126.200 ;
        RECT 163.800 126.100 164.200 126.600 ;
        RECT 163.000 125.800 164.200 126.100 ;
        RECT 164.600 125.800 165.000 126.600 ;
        RECT 165.400 126.500 166.100 126.900 ;
        RECT 166.400 126.800 167.400 127.200 ;
        RECT 169.400 126.800 169.800 127.200 ;
        RECT 171.400 127.100 172.200 127.200 ;
        RECT 173.500 127.100 173.800 128.200 ;
        RECT 178.300 127.700 178.700 127.800 ;
        RECT 179.800 127.700 180.200 129.900 ;
        RECT 178.300 127.400 180.200 127.700 ;
        RECT 175.000 127.100 175.400 127.200 ;
        RECT 176.300 127.100 176.700 127.200 ;
        RECT 171.400 126.800 176.900 127.100 ;
        RECT 165.400 125.500 165.700 126.500 ;
        RECT 163.800 125.200 165.700 125.500 ;
        RECT 166.400 125.200 166.700 126.800 ;
        RECT 167.000 125.400 167.400 126.200 ;
        RECT 168.600 125.400 169.000 126.200 ;
        RECT 161.100 121.100 162.100 125.100 ;
        RECT 163.800 123.500 164.100 125.200 ;
        RECT 166.200 124.900 166.700 125.200 ;
        RECT 169.400 125.100 169.700 126.800 ;
        RECT 172.900 126.700 173.300 126.800 ;
        RECT 172.100 126.200 172.500 126.300 ;
        RECT 173.400 126.200 173.800 126.300 ;
        RECT 176.600 126.200 176.900 126.800 ;
        RECT 177.400 126.400 177.800 126.500 ;
        RECT 172.100 125.900 174.600 126.200 ;
        RECT 174.200 125.800 174.600 125.900 ;
        RECT 176.600 125.800 177.000 126.200 ;
        RECT 177.400 126.100 179.300 126.400 ;
        RECT 178.900 126.000 179.300 126.100 ;
        RECT 171.000 125.500 173.800 125.600 ;
        RECT 171.000 125.400 173.900 125.500 ;
        RECT 171.000 125.300 175.900 125.400 ;
        RECT 165.900 124.600 166.700 124.900 ;
        RECT 168.900 124.700 169.800 125.100 ;
        RECT 163.800 121.500 164.200 123.500 ;
        RECT 165.900 121.100 166.300 124.600 ;
        RECT 168.900 122.200 169.300 124.700 ;
        RECT 168.600 121.800 169.300 122.200 ;
        RECT 168.900 121.100 169.300 121.800 ;
        RECT 171.000 121.100 171.400 125.300 ;
        RECT 173.500 125.100 175.900 125.300 ;
        RECT 172.600 124.500 175.300 124.800 ;
        RECT 172.600 124.400 173.000 124.500 ;
        RECT 174.900 124.400 175.300 124.500 ;
        RECT 175.600 124.500 175.900 125.100 ;
        RECT 176.600 125.200 176.900 125.800 ;
        RECT 178.100 125.700 178.500 125.800 ;
        RECT 179.800 125.700 180.200 127.400 ;
        RECT 178.100 125.400 180.200 125.700 ;
        RECT 176.600 124.900 177.800 125.200 ;
        RECT 176.300 124.500 176.700 124.600 ;
        RECT 175.600 124.200 176.700 124.500 ;
        RECT 177.500 124.400 177.800 124.900 ;
        RECT 177.500 124.000 178.200 124.400 ;
        RECT 174.300 123.700 174.700 123.800 ;
        RECT 175.700 123.700 176.100 123.800 ;
        RECT 172.600 123.100 173.000 123.500 ;
        RECT 174.300 123.400 176.100 123.700 ;
        RECT 175.400 123.100 175.700 123.400 ;
        RECT 177.400 123.100 177.800 123.500 ;
        RECT 172.600 122.800 173.600 123.100 ;
        RECT 173.200 121.100 173.600 122.800 ;
        RECT 175.400 121.100 175.800 123.100 ;
        RECT 177.500 121.100 178.100 123.100 ;
        RECT 179.800 121.100 180.200 125.400 ;
        RECT 2.500 117.200 2.900 119.900 ;
        RECT 4.600 117.500 5.000 119.500 ;
        RECT 2.500 116.800 3.400 117.200 ;
        RECT 2.500 116.400 2.900 116.800 ;
        RECT 2.100 116.100 2.900 116.400 ;
        RECT 1.400 114.800 1.800 115.600 ;
        RECT 2.100 114.200 2.400 116.100 ;
        RECT 4.700 115.800 5.000 117.500 ;
        RECT 3.100 115.500 5.000 115.800 ;
        RECT 3.100 114.500 3.400 115.500 ;
        RECT 1.400 113.800 2.400 114.200 ;
        RECT 2.700 114.100 3.400 114.500 ;
        RECT 3.800 114.400 4.200 115.200 ;
        RECT 4.600 114.400 5.000 115.200 ;
        RECT 5.400 115.100 5.800 119.900 ;
        RECT 7.000 115.700 7.400 119.900 ;
        RECT 9.200 118.200 9.600 119.900 ;
        RECT 8.600 117.900 9.600 118.200 ;
        RECT 11.400 117.900 11.800 119.900 ;
        RECT 13.500 117.900 14.100 119.900 ;
        RECT 8.600 117.500 9.000 117.900 ;
        RECT 11.400 117.600 11.700 117.900 ;
        RECT 10.300 117.300 12.100 117.600 ;
        RECT 13.400 117.500 13.800 117.900 ;
        RECT 10.300 117.200 10.700 117.300 ;
        RECT 11.700 117.200 12.100 117.300 ;
        RECT 8.600 116.500 9.000 116.600 ;
        RECT 10.900 116.500 11.300 116.600 ;
        RECT 8.600 116.200 11.300 116.500 ;
        RECT 11.600 116.500 12.700 116.800 ;
        RECT 11.600 115.900 11.900 116.500 ;
        RECT 12.300 116.400 12.700 116.500 ;
        RECT 13.500 116.600 14.200 117.000 ;
        RECT 13.500 116.100 13.800 116.600 ;
        RECT 9.500 115.700 11.900 115.900 ;
        RECT 7.000 115.600 11.900 115.700 ;
        RECT 12.600 115.800 13.800 116.100 ;
        RECT 7.000 115.500 9.900 115.600 ;
        RECT 7.000 115.400 9.800 115.500 ;
        RECT 12.600 115.200 12.900 115.800 ;
        RECT 15.800 115.600 16.200 119.900 ;
        RECT 16.600 116.200 17.000 119.900 ;
        RECT 18.200 116.200 18.600 119.900 ;
        RECT 16.600 115.900 18.600 116.200 ;
        RECT 19.000 115.900 19.400 119.900 ;
        RECT 20.100 116.300 20.500 119.900 ;
        RECT 20.100 115.900 21.000 116.300 ;
        RECT 14.100 115.300 16.200 115.600 ;
        RECT 14.100 115.200 14.500 115.300 ;
        RECT 6.200 115.100 6.600 115.200 ;
        RECT 10.200 115.100 10.600 115.200 ;
        RECT 5.400 114.800 6.600 115.100 ;
        RECT 8.100 114.800 10.600 115.100 ;
        RECT 12.600 114.800 13.000 115.200 ;
        RECT 14.900 114.900 15.300 115.000 ;
        RECT 2.100 113.500 2.400 113.800 ;
        RECT 2.900 113.900 3.400 114.100 ;
        RECT 2.900 113.600 5.000 113.900 ;
        RECT 2.100 113.300 2.500 113.500 ;
        RECT 2.100 113.000 2.900 113.300 ;
        RECT 2.500 111.500 2.900 113.000 ;
        RECT 4.700 112.500 5.000 113.600 ;
        RECT 4.600 111.500 5.000 112.500 ;
        RECT 5.400 111.100 5.800 114.800 ;
        RECT 8.100 114.700 8.500 114.800 ;
        RECT 9.400 114.700 9.800 114.800 ;
        RECT 8.900 114.200 9.300 114.300 ;
        RECT 12.600 114.200 12.900 114.800 ;
        RECT 13.400 114.600 15.300 114.900 ;
        RECT 13.400 114.500 13.800 114.600 ;
        RECT 7.400 113.900 12.900 114.200 ;
        RECT 7.400 113.800 8.200 113.900 ;
        RECT 6.200 112.400 6.600 113.200 ;
        RECT 7.000 111.100 7.400 113.500 ;
        RECT 9.500 112.800 9.800 113.900 ;
        RECT 12.300 113.800 12.700 113.900 ;
        RECT 15.800 113.600 16.200 115.300 ;
        RECT 17.000 115.200 17.400 115.400 ;
        RECT 19.000 115.200 19.300 115.900 ;
        RECT 16.600 114.900 17.400 115.200 ;
        RECT 18.200 114.900 19.400 115.200 ;
        RECT 16.600 114.800 17.000 114.900 ;
        RECT 17.400 113.800 17.800 114.600 ;
        RECT 14.300 113.300 16.200 113.600 ;
        RECT 14.300 113.200 14.700 113.300 ;
        RECT 8.600 112.100 9.000 112.500 ;
        RECT 9.400 112.400 9.800 112.800 ;
        RECT 10.300 112.700 10.700 112.800 ;
        RECT 10.300 112.400 11.700 112.700 ;
        RECT 11.400 112.100 11.700 112.400 ;
        RECT 13.400 112.100 13.800 112.500 ;
        RECT 8.600 111.800 9.600 112.100 ;
        RECT 9.200 111.100 9.600 111.800 ;
        RECT 11.400 111.100 11.800 112.100 ;
        RECT 13.400 111.800 14.100 112.100 ;
        RECT 13.500 111.100 14.100 111.800 ;
        RECT 15.800 111.100 16.200 113.300 ;
        RECT 18.200 113.100 18.500 114.900 ;
        RECT 19.000 114.800 19.400 114.900 ;
        RECT 19.800 114.800 20.200 115.600 ;
        RECT 20.600 114.200 20.900 115.900 ;
        RECT 22.200 115.700 22.600 119.900 ;
        RECT 24.400 118.200 24.800 119.900 ;
        RECT 23.800 117.900 24.800 118.200 ;
        RECT 26.600 117.900 27.000 119.900 ;
        RECT 28.700 117.900 29.300 119.900 ;
        RECT 23.800 117.500 24.200 117.900 ;
        RECT 26.600 117.600 26.900 117.900 ;
        RECT 25.500 117.300 27.300 117.600 ;
        RECT 28.600 117.500 29.000 117.900 ;
        RECT 25.500 117.200 25.900 117.300 ;
        RECT 26.900 117.200 27.300 117.300 ;
        RECT 23.800 116.500 24.200 116.600 ;
        RECT 26.100 116.500 26.500 116.600 ;
        RECT 23.800 116.200 26.500 116.500 ;
        RECT 26.800 116.500 27.900 116.800 ;
        RECT 26.800 115.900 27.100 116.500 ;
        RECT 27.500 116.400 27.900 116.500 ;
        RECT 28.700 116.600 29.400 117.000 ;
        RECT 28.700 116.100 29.000 116.600 ;
        RECT 24.700 115.700 27.100 115.900 ;
        RECT 22.200 115.600 27.100 115.700 ;
        RECT 27.800 115.800 29.000 116.100 ;
        RECT 22.200 115.500 25.100 115.600 ;
        RECT 22.200 115.400 25.000 115.500 ;
        RECT 25.400 115.100 25.800 115.200 ;
        RECT 23.300 114.800 25.800 115.100 ;
        RECT 27.000 115.100 27.400 115.200 ;
        RECT 27.800 115.100 28.100 115.800 ;
        RECT 31.000 115.600 31.400 119.900 ;
        RECT 31.800 116.200 32.200 119.900 ;
        RECT 33.400 116.200 33.800 119.900 ;
        RECT 31.800 115.900 33.800 116.200 ;
        RECT 34.200 115.900 34.600 119.900 ;
        RECT 35.300 116.300 35.700 119.900 ;
        RECT 35.300 115.900 36.200 116.300 ;
        RECT 29.300 115.300 31.400 115.600 ;
        RECT 29.300 115.200 29.700 115.300 ;
        RECT 27.000 114.800 28.100 115.100 ;
        RECT 30.100 114.900 30.500 115.000 ;
        RECT 23.300 114.700 23.700 114.800 ;
        RECT 24.100 114.200 24.500 114.300 ;
        RECT 27.800 114.200 28.100 114.800 ;
        RECT 28.600 114.600 30.500 114.900 ;
        RECT 28.600 114.500 29.000 114.600 ;
        RECT 20.600 113.800 21.000 114.200 ;
        RECT 22.600 113.900 28.100 114.200 ;
        RECT 22.600 113.800 23.400 113.900 ;
        RECT 19.000 113.100 19.400 113.200 ;
        RECT 20.600 113.100 20.900 113.800 ;
        RECT 18.200 111.100 18.600 113.100 ;
        RECT 19.000 112.800 20.900 113.100 ;
        RECT 18.900 112.400 19.300 112.800 ;
        RECT 20.600 112.100 20.900 112.800 ;
        RECT 21.400 112.400 21.800 113.200 ;
        RECT 20.600 111.100 21.000 112.100 ;
        RECT 22.200 111.100 22.600 113.500 ;
        RECT 24.700 113.200 25.000 113.900 ;
        RECT 27.500 113.800 27.900 113.900 ;
        RECT 31.000 113.600 31.400 115.300 ;
        RECT 32.200 115.200 32.600 115.400 ;
        RECT 34.200 115.200 34.500 115.900 ;
        RECT 31.800 114.900 32.600 115.200 ;
        RECT 33.400 114.900 34.600 115.200 ;
        RECT 31.800 114.800 32.200 114.900 ;
        RECT 32.600 113.800 33.000 114.600 ;
        RECT 29.500 113.300 31.400 113.600 ;
        RECT 29.500 113.200 29.900 113.300 ;
        RECT 23.800 112.100 24.200 112.500 ;
        RECT 24.600 112.400 25.000 113.200 ;
        RECT 25.500 112.700 25.900 112.800 ;
        RECT 25.500 112.400 26.900 112.700 ;
        RECT 26.600 112.100 26.900 112.400 ;
        RECT 28.600 112.100 29.000 112.500 ;
        RECT 23.800 111.800 24.800 112.100 ;
        RECT 24.400 111.100 24.800 111.800 ;
        RECT 26.600 111.100 27.000 112.100 ;
        RECT 28.600 111.800 29.300 112.100 ;
        RECT 28.700 111.100 29.300 111.800 ;
        RECT 31.000 111.100 31.400 113.300 ;
        RECT 33.400 113.200 33.700 114.900 ;
        RECT 34.200 114.800 34.600 114.900 ;
        RECT 35.000 114.800 35.400 115.600 ;
        RECT 35.800 114.200 36.100 115.900 ;
        RECT 35.800 113.800 36.200 114.200 ;
        RECT 36.600 114.100 37.000 114.200 ;
        RECT 39.000 114.100 39.400 114.200 ;
        RECT 36.600 113.800 39.400 114.100 ;
        RECT 33.400 111.100 33.800 113.200 ;
        RECT 34.200 113.100 34.600 113.200 ;
        RECT 35.800 113.100 36.100 113.800 ;
        RECT 39.000 113.400 39.400 113.800 ;
        RECT 34.200 112.800 36.100 113.100 ;
        RECT 34.100 112.400 34.500 112.800 ;
        RECT 35.800 112.100 36.100 112.800 ;
        RECT 36.600 112.400 37.000 113.200 ;
        RECT 39.800 113.100 40.200 119.900 ;
        RECT 41.400 117.500 41.800 119.500 ;
        RECT 40.600 115.800 41.000 116.600 ;
        RECT 41.400 115.800 41.700 117.500 ;
        RECT 43.500 117.200 43.900 119.900 ;
        RECT 43.500 116.800 44.200 117.200 ;
        RECT 43.500 116.400 43.900 116.800 ;
        RECT 43.500 116.100 44.300 116.400 ;
        RECT 41.400 115.500 43.300 115.800 ;
        RECT 41.400 114.400 41.800 115.200 ;
        RECT 42.200 114.400 42.600 115.200 ;
        RECT 43.000 114.500 43.300 115.500 ;
        RECT 43.000 114.100 43.700 114.500 ;
        RECT 44.000 114.200 44.300 116.100 ;
        RECT 44.600 115.100 45.000 115.600 ;
        RECT 46.200 115.100 46.600 119.900 ;
        RECT 47.800 115.700 48.200 119.900 ;
        RECT 50.000 118.200 50.400 119.900 ;
        RECT 49.400 117.900 50.400 118.200 ;
        RECT 52.200 117.900 52.600 119.900 ;
        RECT 54.300 117.900 54.900 119.900 ;
        RECT 49.400 117.500 49.800 117.900 ;
        RECT 52.200 117.600 52.500 117.900 ;
        RECT 51.100 117.300 52.900 117.600 ;
        RECT 54.200 117.500 54.600 117.900 ;
        RECT 51.100 117.200 51.500 117.300 ;
        RECT 52.500 117.200 52.900 117.300 ;
        RECT 49.400 116.500 49.800 116.600 ;
        RECT 51.700 116.500 52.100 116.600 ;
        RECT 49.400 116.200 52.100 116.500 ;
        RECT 52.400 116.500 53.500 116.800 ;
        RECT 52.400 115.900 52.700 116.500 ;
        RECT 53.100 116.400 53.500 116.500 ;
        RECT 54.300 116.600 55.000 117.000 ;
        RECT 54.300 116.100 54.600 116.600 ;
        RECT 50.300 115.700 52.700 115.900 ;
        RECT 47.800 115.600 52.700 115.700 ;
        RECT 53.400 115.800 54.600 116.100 ;
        RECT 47.800 115.500 50.700 115.600 ;
        RECT 47.800 115.400 50.600 115.500 ;
        RECT 51.000 115.100 51.400 115.200 ;
        RECT 44.600 114.800 46.600 115.100 ;
        RECT 43.000 113.900 43.500 114.100 ;
        RECT 41.400 113.600 43.500 113.900 ;
        RECT 44.000 113.800 45.000 114.200 ;
        RECT 39.800 112.800 40.700 113.100 ;
        RECT 35.800 111.100 36.200 112.100 ;
        RECT 40.300 111.100 40.700 112.800 ;
        RECT 41.400 112.500 41.700 113.600 ;
        RECT 44.000 113.500 44.300 113.800 ;
        RECT 43.900 113.300 44.300 113.500 ;
        RECT 43.500 113.000 44.300 113.300 ;
        RECT 41.400 111.500 41.800 112.500 ;
        RECT 43.500 111.500 43.900 113.000 ;
        RECT 46.200 111.100 46.600 114.800 ;
        RECT 48.900 114.800 51.400 115.100 ;
        RECT 48.900 114.700 49.300 114.800 ;
        RECT 50.200 114.700 50.600 114.800 ;
        RECT 49.700 114.200 50.100 114.300 ;
        RECT 53.400 114.200 53.700 115.800 ;
        RECT 55.000 115.600 55.400 116.200 ;
        RECT 56.600 115.600 57.000 119.900 ;
        RECT 54.900 115.300 57.000 115.600 ;
        RECT 54.900 115.200 55.300 115.300 ;
        RECT 55.700 114.900 56.100 115.000 ;
        RECT 54.200 114.600 56.100 114.900 ;
        RECT 54.200 114.500 54.600 114.600 ;
        RECT 48.200 113.900 53.700 114.200 ;
        RECT 48.200 113.800 49.000 113.900 ;
        RECT 47.000 112.400 47.400 113.200 ;
        RECT 47.800 111.100 48.200 113.500 ;
        RECT 50.300 112.800 50.600 113.900 ;
        RECT 51.000 113.800 51.400 113.900 ;
        RECT 53.100 113.800 53.500 113.900 ;
        RECT 56.600 113.600 57.000 115.300 ;
        RECT 55.100 113.300 57.000 113.600 ;
        RECT 55.100 113.200 55.500 113.300 ;
        RECT 49.400 112.100 49.800 112.500 ;
        RECT 50.200 112.400 50.600 112.800 ;
        RECT 51.100 112.700 51.500 112.800 ;
        RECT 51.100 112.400 52.500 112.700 ;
        RECT 52.200 112.100 52.500 112.400 ;
        RECT 54.200 112.100 54.600 112.500 ;
        RECT 49.400 111.800 50.400 112.100 ;
        RECT 50.000 111.100 50.400 111.800 ;
        RECT 52.200 111.100 52.600 112.100 ;
        RECT 54.200 111.800 54.900 112.100 ;
        RECT 54.300 111.100 54.900 111.800 ;
        RECT 56.600 111.100 57.000 113.300 ;
        RECT 57.400 115.600 57.800 119.900 ;
        RECT 59.500 117.900 60.100 119.900 ;
        RECT 61.800 117.900 62.200 119.900 ;
        RECT 64.000 118.200 64.400 119.900 ;
        RECT 64.000 117.900 65.000 118.200 ;
        RECT 59.800 117.500 60.200 117.900 ;
        RECT 61.900 117.600 62.200 117.900 ;
        RECT 61.500 117.300 63.300 117.600 ;
        RECT 64.600 117.500 65.000 117.900 ;
        RECT 61.500 117.200 61.900 117.300 ;
        RECT 62.900 117.200 63.300 117.300 ;
        RECT 59.400 116.600 60.100 117.000 ;
        RECT 59.800 116.100 60.100 116.600 ;
        RECT 60.900 116.500 62.000 116.800 ;
        RECT 60.900 116.400 61.300 116.500 ;
        RECT 59.800 115.800 61.000 116.100 ;
        RECT 57.400 115.300 59.500 115.600 ;
        RECT 57.400 113.600 57.800 115.300 ;
        RECT 59.100 115.200 59.500 115.300 ;
        RECT 58.300 114.900 58.700 115.000 ;
        RECT 58.300 114.600 60.200 114.900 ;
        RECT 59.800 114.500 60.200 114.600 ;
        RECT 60.700 114.200 61.000 115.800 ;
        RECT 61.700 115.900 62.000 116.500 ;
        RECT 62.300 116.500 62.700 116.600 ;
        RECT 64.600 116.500 65.000 116.600 ;
        RECT 62.300 116.200 65.000 116.500 ;
        RECT 61.700 115.700 64.100 115.900 ;
        RECT 66.200 115.700 66.600 119.900 ;
        RECT 61.700 115.600 66.600 115.700 ;
        RECT 63.700 115.500 66.600 115.600 ;
        RECT 63.800 115.400 66.600 115.500 ;
        RECT 63.000 115.100 63.400 115.200 ;
        RECT 67.800 115.100 68.200 119.900 ;
        RECT 70.500 116.400 70.900 119.900 ;
        RECT 72.600 117.500 73.000 119.500 ;
        RECT 70.100 116.100 70.900 116.400 ;
        RECT 69.400 115.100 69.800 115.600 ;
        RECT 63.000 114.800 65.500 115.100 ;
        RECT 65.100 114.700 65.500 114.800 ;
        RECT 67.800 114.800 69.800 115.100 ;
        RECT 64.300 114.200 64.700 114.300 ;
        RECT 60.700 113.900 66.200 114.200 ;
        RECT 60.900 113.800 61.300 113.900 ;
        RECT 57.400 113.300 59.300 113.600 ;
        RECT 57.400 111.100 57.800 113.300 ;
        RECT 58.900 113.200 59.300 113.300 ;
        RECT 63.800 112.800 64.100 113.900 ;
        RECT 65.400 113.800 66.200 113.900 ;
        RECT 62.900 112.700 63.300 112.800 ;
        RECT 59.800 112.100 60.200 112.500 ;
        RECT 61.900 112.400 63.300 112.700 ;
        RECT 63.800 112.400 64.200 112.800 ;
        RECT 61.900 112.100 62.200 112.400 ;
        RECT 64.600 112.100 65.000 112.500 ;
        RECT 59.500 111.800 60.200 112.100 ;
        RECT 59.500 111.100 60.100 111.800 ;
        RECT 61.800 111.100 62.200 112.100 ;
        RECT 64.000 111.800 65.000 112.100 ;
        RECT 64.000 111.100 64.400 111.800 ;
        RECT 66.200 111.100 66.600 113.500 ;
        RECT 67.000 112.400 67.400 113.200 ;
        RECT 67.800 111.100 68.200 114.800 ;
        RECT 70.100 114.200 70.400 116.100 ;
        RECT 72.700 115.800 73.000 117.500 ;
        RECT 73.400 116.900 73.800 119.900 ;
        RECT 73.500 116.600 73.800 116.900 ;
        RECT 75.000 119.600 77.000 119.900 ;
        RECT 75.000 116.900 75.400 119.600 ;
        RECT 75.800 116.900 76.200 119.300 ;
        RECT 76.600 117.000 77.000 119.600 ;
        RECT 77.500 119.600 79.300 119.900 ;
        RECT 77.500 119.500 77.800 119.600 ;
        RECT 75.000 116.600 75.300 116.900 ;
        RECT 73.500 116.300 75.300 116.600 ;
        RECT 75.900 116.700 76.200 116.900 ;
        RECT 77.400 116.700 77.800 119.500 ;
        RECT 79.000 119.500 79.300 119.600 ;
        RECT 75.900 116.500 77.800 116.700 ;
        RECT 78.200 116.500 78.600 119.300 ;
        RECT 79.000 116.500 79.400 119.500 ;
        RECT 79.800 117.900 80.200 119.900 ;
        RECT 79.900 117.800 80.200 117.900 ;
        RECT 81.400 117.900 81.800 119.900 ;
        RECT 81.400 117.800 81.700 117.900 ;
        RECT 79.900 117.500 81.700 117.800 ;
        RECT 75.900 116.400 77.700 116.500 ;
        RECT 78.200 116.200 78.500 116.500 ;
        RECT 79.900 116.200 80.200 117.500 ;
        RECT 80.600 116.400 81.000 117.200 ;
        RECT 78.200 116.100 78.600 116.200 ;
        RECT 71.100 115.500 73.000 115.800 ;
        RECT 76.900 115.800 78.600 116.100 ;
        RECT 79.800 115.800 80.200 116.200 ;
        RECT 81.400 116.100 81.800 116.200 ;
        RECT 82.200 116.100 82.600 116.200 ;
        RECT 81.400 115.800 82.600 116.100 ;
        RECT 83.000 115.800 83.400 116.600 ;
        RECT 71.100 114.500 71.400 115.500 ;
        RECT 69.400 113.800 70.400 114.200 ;
        RECT 70.700 114.100 71.400 114.500 ;
        RECT 71.800 114.400 72.200 115.200 ;
        RECT 72.600 114.400 73.000 115.200 ;
        RECT 75.800 114.800 76.600 115.200 ;
        RECT 70.100 113.500 70.400 113.800 ;
        RECT 70.900 113.900 71.400 114.100 ;
        RECT 73.400 114.100 73.800 114.200 ;
        RECT 75.000 114.100 75.800 114.200 ;
        RECT 70.900 113.600 73.000 113.900 ;
        RECT 73.400 113.800 75.800 114.100 ;
        RECT 70.100 113.300 70.500 113.500 ;
        RECT 70.100 113.000 70.900 113.300 ;
        RECT 70.500 112.200 70.900 113.000 ;
        RECT 72.700 112.500 73.000 113.600 ;
        RECT 74.200 112.800 75.100 113.200 ;
        RECT 76.900 112.500 77.200 115.800 ;
        RECT 79.900 114.200 80.200 115.800 ;
        RECT 82.200 115.400 82.600 115.800 ;
        RECT 81.000 114.800 81.800 115.200 ;
        RECT 79.900 114.100 80.700 114.200 ;
        RECT 79.900 113.900 80.800 114.100 ;
        RECT 70.500 111.800 71.400 112.200 ;
        RECT 70.500 111.500 70.900 111.800 ;
        RECT 72.600 111.500 73.000 112.500 ;
        RECT 75.200 112.200 77.200 112.500 ;
        RECT 75.200 112.100 75.500 112.200 ;
        RECT 75.000 111.800 75.500 112.100 ;
        RECT 76.600 112.100 77.200 112.200 ;
        RECT 79.000 112.100 79.400 112.200 ;
        RECT 76.600 111.800 79.400 112.100 ;
        RECT 75.000 111.100 75.400 111.800 ;
        RECT 76.600 111.100 77.000 111.800 ;
        RECT 80.400 111.100 80.800 113.900 ;
        RECT 83.000 113.800 83.400 114.200 ;
        RECT 83.000 113.200 83.300 113.800 ;
        RECT 83.800 113.200 84.200 119.900 ;
        RECT 85.400 117.500 85.800 119.500 ;
        RECT 85.400 115.800 85.700 117.500 ;
        RECT 87.500 116.400 87.900 119.900 ;
        RECT 87.500 116.100 88.300 116.400 ;
        RECT 85.400 115.500 87.300 115.800 ;
        RECT 85.400 114.400 85.800 115.200 ;
        RECT 86.200 114.400 86.600 115.200 ;
        RECT 87.000 114.500 87.300 115.500 ;
        RECT 84.600 113.400 85.000 114.200 ;
        RECT 87.000 114.100 87.700 114.500 ;
        RECT 88.000 114.200 88.300 116.100 ;
        RECT 88.600 115.100 89.000 115.600 ;
        RECT 91.800 115.100 92.200 119.900 ;
        RECT 93.400 116.200 93.800 119.900 ;
        RECT 95.000 119.600 97.000 119.900 ;
        RECT 95.000 116.200 95.400 119.600 ;
        RECT 93.400 115.900 95.400 116.200 ;
        RECT 95.800 115.900 96.200 119.300 ;
        RECT 96.600 115.900 97.000 119.600 ;
        RECT 95.800 115.600 96.100 115.900 ;
        RECT 97.400 115.800 97.800 116.600 ;
        RECT 93.800 115.200 94.200 115.400 ;
        RECT 95.100 115.300 96.100 115.600 ;
        RECT 95.100 115.200 95.400 115.300 ;
        RECT 88.600 114.800 92.200 115.100 ;
        RECT 92.600 115.100 93.000 115.200 ;
        RECT 93.400 115.100 94.200 115.200 ;
        RECT 92.600 114.900 94.200 115.100 ;
        RECT 92.600 114.800 93.800 114.900 ;
        RECT 95.000 114.800 95.400 115.200 ;
        RECT 96.600 114.800 97.000 115.600 ;
        RECT 88.000 114.100 89.000 114.200 ;
        RECT 91.000 114.100 91.400 114.200 ;
        RECT 87.000 113.900 87.500 114.100 ;
        RECT 85.400 113.600 87.500 113.900 ;
        RECT 88.000 113.800 91.400 114.100 ;
        RECT 83.000 112.800 84.200 113.200 ;
        RECT 83.300 111.100 83.700 112.800 ;
        RECT 85.400 112.500 85.700 113.600 ;
        RECT 88.000 113.500 88.300 113.800 ;
        RECT 87.900 113.300 88.300 113.500 ;
        RECT 87.500 113.000 88.300 113.300 ;
        RECT 85.400 111.500 85.800 112.500 ;
        RECT 87.500 111.500 87.900 113.000 ;
        RECT 91.800 111.100 92.200 114.800 ;
        RECT 93.400 114.100 93.800 114.200 ;
        RECT 94.200 114.100 94.600 114.600 ;
        RECT 93.400 113.800 94.600 114.100 ;
        RECT 92.600 112.400 93.000 113.200 ;
        RECT 95.100 113.100 95.400 114.800 ;
        RECT 95.700 114.400 96.100 114.800 ;
        RECT 95.800 114.200 96.100 114.400 ;
        RECT 95.800 113.800 96.200 114.200 ;
        RECT 98.200 113.100 98.600 119.900 ;
        RECT 99.800 115.600 100.200 119.900 ;
        RECT 101.900 117.900 102.500 119.900 ;
        RECT 104.200 117.900 104.600 119.900 ;
        RECT 106.400 118.200 106.800 119.900 ;
        RECT 106.400 117.900 107.400 118.200 ;
        RECT 102.200 117.500 102.600 117.900 ;
        RECT 104.300 117.600 104.600 117.900 ;
        RECT 103.900 117.300 105.700 117.600 ;
        RECT 107.000 117.500 107.400 117.900 ;
        RECT 103.900 117.200 104.300 117.300 ;
        RECT 105.300 117.200 105.700 117.300 ;
        RECT 101.800 116.600 102.500 117.000 ;
        RECT 102.200 116.100 102.500 116.600 ;
        RECT 103.300 116.500 104.400 116.800 ;
        RECT 103.300 116.400 103.700 116.500 ;
        RECT 102.200 115.800 103.400 116.100 ;
        RECT 99.800 115.300 101.900 115.600 ;
        RECT 99.000 113.400 99.400 114.200 ;
        RECT 99.800 113.600 100.200 115.300 ;
        RECT 101.500 115.200 101.900 115.300 ;
        RECT 100.700 114.900 101.100 115.000 ;
        RECT 100.700 114.600 102.600 114.900 ;
        RECT 102.200 114.500 102.600 114.600 ;
        RECT 103.100 114.200 103.400 115.800 ;
        RECT 104.100 115.900 104.400 116.500 ;
        RECT 104.700 116.500 105.100 116.600 ;
        RECT 107.000 116.500 107.400 116.600 ;
        RECT 104.700 116.200 107.400 116.500 ;
        RECT 104.100 115.700 106.500 115.900 ;
        RECT 108.600 115.700 109.000 119.900 ;
        RECT 104.100 115.600 109.000 115.700 ;
        RECT 106.100 115.500 109.000 115.600 ;
        RECT 106.200 115.400 109.000 115.500 ;
        RECT 105.400 115.100 105.800 115.200 ;
        RECT 110.200 115.100 110.600 119.900 ;
        RECT 112.900 116.400 113.300 119.900 ;
        RECT 115.000 117.500 115.400 119.500 ;
        RECT 112.500 116.100 113.300 116.400 ;
        RECT 112.500 115.800 113.000 116.100 ;
        RECT 115.100 115.800 115.400 117.500 ;
        RECT 111.800 115.100 112.200 115.600 ;
        RECT 105.400 114.800 107.900 115.100 ;
        RECT 107.500 114.700 107.900 114.800 ;
        RECT 110.200 114.800 112.200 115.100 ;
        RECT 106.700 114.200 107.100 114.300 ;
        RECT 103.100 113.900 108.600 114.200 ;
        RECT 103.300 113.800 103.700 113.900 ;
        RECT 105.400 113.800 105.800 113.900 ;
        RECT 94.900 111.100 95.700 113.100 ;
        RECT 97.700 112.800 98.600 113.100 ;
        RECT 99.800 113.300 101.700 113.600 ;
        RECT 97.700 112.200 98.100 112.800 ;
        RECT 97.400 111.800 98.100 112.200 ;
        RECT 97.700 111.100 98.100 111.800 ;
        RECT 99.800 111.100 100.200 113.300 ;
        RECT 101.300 113.200 101.700 113.300 ;
        RECT 106.200 112.800 106.500 113.900 ;
        RECT 107.800 113.800 108.600 113.900 ;
        RECT 105.300 112.700 105.700 112.800 ;
        RECT 102.200 112.100 102.600 112.500 ;
        RECT 104.300 112.400 105.700 112.700 ;
        RECT 106.200 112.400 106.600 112.800 ;
        RECT 104.300 112.100 104.600 112.400 ;
        RECT 107.000 112.100 107.400 112.500 ;
        RECT 101.900 111.800 102.600 112.100 ;
        RECT 101.900 111.100 102.500 111.800 ;
        RECT 104.200 111.100 104.600 112.100 ;
        RECT 106.400 111.800 107.400 112.100 ;
        RECT 106.400 111.100 106.800 111.800 ;
        RECT 108.600 111.100 109.000 113.500 ;
        RECT 109.400 112.400 109.800 113.200 ;
        RECT 110.200 111.100 110.600 114.800 ;
        RECT 112.500 114.200 112.800 115.800 ;
        RECT 113.500 115.500 115.400 115.800 ;
        RECT 115.800 115.600 116.200 119.900 ;
        RECT 117.900 117.900 118.500 119.900 ;
        RECT 120.200 117.900 120.600 119.900 ;
        RECT 122.400 118.200 122.800 119.900 ;
        RECT 122.400 117.900 123.400 118.200 ;
        RECT 118.200 117.500 118.600 117.900 ;
        RECT 120.300 117.600 120.600 117.900 ;
        RECT 119.900 117.300 121.700 117.600 ;
        RECT 123.000 117.500 123.400 117.900 ;
        RECT 119.900 117.200 120.300 117.300 ;
        RECT 121.300 117.200 121.700 117.300 ;
        RECT 117.800 116.600 118.500 117.000 ;
        RECT 118.200 116.100 118.500 116.600 ;
        RECT 119.300 116.500 120.400 116.800 ;
        RECT 119.300 116.400 119.700 116.500 ;
        RECT 118.200 115.800 119.400 116.100 ;
        RECT 113.500 114.500 113.800 115.500 ;
        RECT 115.800 115.300 117.900 115.600 ;
        RECT 111.800 113.800 112.800 114.200 ;
        RECT 113.100 114.100 113.800 114.500 ;
        RECT 114.200 114.400 114.600 115.200 ;
        RECT 115.000 114.400 115.400 115.200 ;
        RECT 112.500 113.500 112.800 113.800 ;
        RECT 113.300 113.900 113.800 114.100 ;
        RECT 113.300 113.600 115.400 113.900 ;
        RECT 112.500 113.300 112.900 113.500 ;
        RECT 112.500 113.000 113.300 113.300 ;
        RECT 112.900 111.500 113.300 113.000 ;
        RECT 115.100 112.500 115.400 113.600 ;
        RECT 115.000 111.500 115.400 112.500 ;
        RECT 115.800 113.600 116.200 115.300 ;
        RECT 117.500 115.200 117.900 115.300 ;
        RECT 116.700 114.900 117.100 115.000 ;
        RECT 116.700 114.600 118.600 114.900 ;
        RECT 118.200 114.500 118.600 114.600 ;
        RECT 119.100 114.200 119.400 115.800 ;
        RECT 120.100 115.900 120.400 116.500 ;
        RECT 120.700 116.500 121.100 116.600 ;
        RECT 123.000 116.500 123.400 116.600 ;
        RECT 120.700 116.200 123.400 116.500 ;
        RECT 120.100 115.700 122.500 115.900 ;
        RECT 124.600 115.700 125.000 119.900 ;
        RECT 120.100 115.600 125.000 115.700 ;
        RECT 126.200 115.600 126.600 119.900 ;
        RECT 127.800 115.600 128.200 119.900 ;
        RECT 129.400 115.600 129.800 119.900 ;
        RECT 131.000 115.600 131.400 119.900 ;
        RECT 122.100 115.500 125.000 115.600 ;
        RECT 122.200 115.400 125.000 115.500 ;
        RECT 125.400 115.200 126.600 115.600 ;
        RECT 127.100 115.200 128.200 115.600 ;
        RECT 128.700 115.200 129.800 115.600 ;
        RECT 130.500 115.200 131.400 115.600 ;
        RECT 132.600 117.500 133.000 119.500 ;
        RECT 132.600 115.800 132.900 117.500 ;
        RECT 134.700 116.400 135.100 119.900 ;
        RECT 137.400 117.100 137.800 119.900 ;
        RECT 139.000 117.100 139.400 117.200 ;
        RECT 137.400 116.800 139.400 117.100 ;
        RECT 134.700 116.100 135.500 116.400 ;
        RECT 132.600 115.500 134.500 115.800 ;
        RECT 121.400 115.100 121.800 115.200 ;
        RECT 121.400 114.800 123.900 115.100 ;
        RECT 123.500 114.700 123.900 114.800 ;
        RECT 122.700 114.200 123.100 114.300 ;
        RECT 119.100 113.900 124.600 114.200 ;
        RECT 119.300 113.800 119.700 113.900 ;
        RECT 121.400 113.800 121.800 113.900 ;
        RECT 115.800 113.300 117.700 113.600 ;
        RECT 115.800 111.100 116.200 113.300 ;
        RECT 117.300 113.200 117.700 113.300 ;
        RECT 122.200 112.800 122.500 113.900 ;
        RECT 123.800 113.800 124.600 113.900 ;
        RECT 125.400 113.800 125.800 115.200 ;
        RECT 127.100 114.500 127.500 115.200 ;
        RECT 128.700 114.500 129.100 115.200 ;
        RECT 130.500 114.500 130.900 115.200 ;
        RECT 126.200 114.100 127.500 114.500 ;
        RECT 127.900 114.100 129.100 114.500 ;
        RECT 129.600 114.100 130.900 114.500 ;
        RECT 132.600 114.400 133.000 115.200 ;
        RECT 133.400 114.400 133.800 115.200 ;
        RECT 134.200 114.500 134.500 115.500 ;
        RECT 127.100 113.800 127.500 114.100 ;
        RECT 128.700 113.800 129.100 114.100 ;
        RECT 130.500 113.800 130.900 114.100 ;
        RECT 134.200 114.100 134.900 114.500 ;
        RECT 135.200 114.200 135.500 116.100 ;
        RECT 135.800 115.100 136.200 115.600 ;
        RECT 137.400 115.100 137.800 116.800 ;
        RECT 135.800 114.800 137.800 115.100 ;
        RECT 135.200 114.100 136.200 114.200 ;
        RECT 136.600 114.100 137.000 114.200 ;
        RECT 134.200 113.900 134.700 114.100 ;
        RECT 121.300 112.700 121.700 112.800 ;
        RECT 118.200 112.100 118.600 112.500 ;
        RECT 120.300 112.400 121.700 112.700 ;
        RECT 122.200 112.400 122.600 112.800 ;
        RECT 120.300 112.100 120.600 112.400 ;
        RECT 123.000 112.100 123.400 112.500 ;
        RECT 117.900 111.800 118.600 112.100 ;
        RECT 117.900 111.100 118.500 111.800 ;
        RECT 120.200 111.100 120.600 112.100 ;
        RECT 122.400 111.800 123.400 112.100 ;
        RECT 122.400 111.100 122.800 111.800 ;
        RECT 124.600 111.100 125.000 113.500 ;
        RECT 125.400 113.400 126.600 113.800 ;
        RECT 127.100 113.400 128.200 113.800 ;
        RECT 128.700 113.400 129.800 113.800 ;
        RECT 130.500 113.400 131.400 113.800 ;
        RECT 126.200 111.100 126.600 113.400 ;
        RECT 127.800 111.100 128.200 113.400 ;
        RECT 129.400 111.100 129.800 113.400 ;
        RECT 131.000 111.100 131.400 113.400 ;
        RECT 132.600 113.600 134.700 113.900 ;
        RECT 135.200 113.800 137.000 114.100 ;
        RECT 132.600 112.500 132.900 113.600 ;
        RECT 135.200 113.500 135.500 113.800 ;
        RECT 135.100 113.300 135.500 113.500 ;
        RECT 134.700 113.000 135.500 113.300 ;
        RECT 132.600 111.500 133.000 112.500 ;
        RECT 134.700 111.500 135.100 113.000 ;
        RECT 137.400 111.100 137.800 114.800 ;
        RECT 140.600 115.600 141.000 119.900 ;
        RECT 142.700 117.900 143.300 119.900 ;
        RECT 145.000 117.900 145.400 119.900 ;
        RECT 147.200 118.200 147.600 119.900 ;
        RECT 147.200 117.900 148.200 118.200 ;
        RECT 143.000 117.500 143.400 117.900 ;
        RECT 145.100 117.600 145.400 117.900 ;
        RECT 144.700 117.300 146.500 117.600 ;
        RECT 147.800 117.500 148.200 117.900 ;
        RECT 144.700 117.200 145.100 117.300 ;
        RECT 146.100 117.200 146.500 117.300 ;
        RECT 142.600 116.600 143.300 117.000 ;
        RECT 143.000 116.100 143.300 116.600 ;
        RECT 144.100 116.500 145.200 116.800 ;
        RECT 144.100 116.400 144.500 116.500 ;
        RECT 143.000 115.800 144.200 116.100 ;
        RECT 140.600 115.300 142.700 115.600 ;
        RECT 140.600 113.600 141.000 115.300 ;
        RECT 142.300 115.200 142.700 115.300 ;
        RECT 143.900 115.200 144.200 115.800 ;
        RECT 144.900 115.900 145.200 116.500 ;
        RECT 145.500 116.500 145.900 116.600 ;
        RECT 147.800 116.500 148.200 116.600 ;
        RECT 145.500 116.200 148.200 116.500 ;
        RECT 144.900 115.700 147.300 115.900 ;
        RECT 149.400 115.700 149.800 119.900 ;
        RECT 144.900 115.600 149.800 115.700 ;
        RECT 146.900 115.500 149.800 115.600 ;
        RECT 147.000 115.400 149.800 115.500 ;
        RECT 141.500 114.900 141.900 115.000 ;
        RECT 141.500 114.600 143.400 114.900 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 146.200 115.100 146.600 115.200 ;
        RECT 146.200 114.800 148.700 115.100 ;
        RECT 143.000 114.500 143.400 114.600 ;
        RECT 143.900 114.200 144.200 114.800 ;
        RECT 148.300 114.700 148.700 114.800 ;
        RECT 147.500 114.200 147.900 114.300 ;
        RECT 143.900 113.900 149.400 114.200 ;
        RECT 144.100 113.800 144.500 113.900 ;
        RECT 140.600 113.300 142.500 113.600 ;
        RECT 138.200 113.100 138.600 113.200 ;
        RECT 138.200 112.800 140.100 113.100 ;
        RECT 138.200 112.400 138.600 112.800 ;
        RECT 139.800 112.100 140.100 112.800 ;
        RECT 140.600 112.100 141.000 113.300 ;
        RECT 142.100 113.200 142.500 113.300 ;
        RECT 147.000 112.800 147.300 113.900 ;
        RECT 148.600 113.800 149.400 113.900 ;
        RECT 146.100 112.700 146.500 112.800 ;
        RECT 143.000 112.100 143.400 112.500 ;
        RECT 145.100 112.400 146.500 112.700 ;
        RECT 147.000 112.400 147.400 112.800 ;
        RECT 145.100 112.100 145.400 112.400 ;
        RECT 147.800 112.100 148.200 112.500 ;
        RECT 139.800 111.800 141.000 112.100 ;
        RECT 140.600 111.100 141.000 111.800 ;
        RECT 142.700 111.800 143.400 112.100 ;
        RECT 142.700 111.100 143.300 111.800 ;
        RECT 145.000 111.100 145.400 112.100 ;
        RECT 147.200 111.800 148.200 112.100 ;
        RECT 147.200 111.100 147.600 111.800 ;
        RECT 149.400 111.100 149.800 113.500 ;
        RECT 150.200 111.100 150.600 119.900 ;
        RECT 151.800 115.700 152.200 119.900 ;
        RECT 154.000 118.200 154.400 119.900 ;
        RECT 153.400 117.900 154.400 118.200 ;
        RECT 156.200 117.900 156.600 119.900 ;
        RECT 158.300 117.900 158.900 119.900 ;
        RECT 153.400 117.500 153.800 117.900 ;
        RECT 156.200 117.600 156.500 117.900 ;
        RECT 155.100 117.300 156.900 117.600 ;
        RECT 158.200 117.500 158.600 117.900 ;
        RECT 155.100 117.200 155.500 117.300 ;
        RECT 156.500 117.200 156.900 117.300 ;
        RECT 153.400 116.500 153.800 116.600 ;
        RECT 155.700 116.500 156.100 116.600 ;
        RECT 153.400 116.200 156.100 116.500 ;
        RECT 156.400 116.500 157.500 116.800 ;
        RECT 156.400 115.900 156.700 116.500 ;
        RECT 157.100 116.400 157.500 116.500 ;
        RECT 158.300 116.600 159.000 117.000 ;
        RECT 158.300 116.100 158.600 116.600 ;
        RECT 154.300 115.700 156.700 115.900 ;
        RECT 151.800 115.600 156.700 115.700 ;
        RECT 157.400 115.800 158.600 116.100 ;
        RECT 151.800 115.500 154.700 115.600 ;
        RECT 151.800 115.400 154.600 115.500 ;
        RECT 155.000 115.100 155.400 115.200 ;
        RECT 152.900 114.800 155.400 115.100 ;
        RECT 152.900 114.700 153.300 114.800 ;
        RECT 153.700 114.200 154.100 114.300 ;
        RECT 157.400 114.200 157.700 115.800 ;
        RECT 160.600 115.600 161.000 119.900 ;
        RECT 158.900 115.300 161.000 115.600 ;
        RECT 161.400 117.500 161.800 119.500 ;
        RECT 161.400 115.800 161.700 117.500 ;
        RECT 163.500 116.400 163.900 119.900 ;
        RECT 163.500 116.100 164.300 116.400 ;
        RECT 161.400 115.500 163.300 115.800 ;
        RECT 158.900 115.200 159.300 115.300 ;
        RECT 159.700 114.900 160.100 115.000 ;
        RECT 158.200 114.600 160.100 114.900 ;
        RECT 158.200 114.500 158.600 114.600 ;
        RECT 152.200 113.900 157.700 114.200 ;
        RECT 152.200 113.800 153.000 113.900 ;
        RECT 151.000 112.400 151.400 113.200 ;
        RECT 151.800 111.100 152.200 113.500 ;
        RECT 154.300 112.800 154.600 113.900 ;
        RECT 157.100 113.800 157.500 113.900 ;
        RECT 160.600 113.600 161.000 115.300 ;
        RECT 161.400 114.400 161.800 115.200 ;
        RECT 162.200 114.400 162.600 115.200 ;
        RECT 163.000 114.500 163.300 115.500 ;
        RECT 163.000 114.100 163.700 114.500 ;
        RECT 164.000 114.200 164.300 116.100 ;
        RECT 164.600 115.100 165.000 115.600 ;
        RECT 166.200 115.100 166.600 119.900 ;
        RECT 164.600 114.800 166.600 115.100 ;
        RECT 163.000 113.900 163.500 114.100 ;
        RECT 159.100 113.300 161.000 113.600 ;
        RECT 159.100 113.200 159.500 113.300 ;
        RECT 153.400 112.100 153.800 112.500 ;
        RECT 154.200 112.400 154.600 112.800 ;
        RECT 155.100 112.700 155.500 112.800 ;
        RECT 155.100 112.400 156.500 112.700 ;
        RECT 156.200 112.100 156.500 112.400 ;
        RECT 158.200 112.100 158.600 112.500 ;
        RECT 153.400 111.800 154.400 112.100 ;
        RECT 154.000 111.100 154.400 111.800 ;
        RECT 156.200 111.100 156.600 112.100 ;
        RECT 158.200 111.800 158.900 112.100 ;
        RECT 158.300 111.100 158.900 111.800 ;
        RECT 160.600 111.100 161.000 113.300 ;
        RECT 161.400 113.600 163.500 113.900 ;
        RECT 164.000 113.800 165.000 114.200 ;
        RECT 161.400 112.500 161.700 113.600 ;
        RECT 164.000 113.500 164.300 113.800 ;
        RECT 163.900 113.300 164.300 113.500 ;
        RECT 163.500 113.200 164.300 113.300 ;
        RECT 163.000 113.000 164.300 113.200 ;
        RECT 163.000 112.800 163.900 113.000 ;
        RECT 161.400 111.500 161.800 112.500 ;
        RECT 163.500 111.500 163.900 112.800 ;
        RECT 166.200 111.100 166.600 114.800 ;
        RECT 167.000 114.100 167.400 114.200 ;
        RECT 167.800 114.100 168.200 114.200 ;
        RECT 167.000 113.800 168.200 114.100 ;
        RECT 167.000 113.200 167.300 113.800 ;
        RECT 167.800 113.400 168.200 113.800 ;
        RECT 167.000 112.400 167.400 113.200 ;
        RECT 168.600 113.100 169.000 119.900 ;
        RECT 169.400 115.800 169.800 116.600 ;
        RECT 171.500 116.200 171.900 119.900 ;
        RECT 172.200 116.800 172.600 117.200 ;
        RECT 173.400 116.900 173.800 119.900 ;
        RECT 172.300 116.200 172.600 116.800 ;
        RECT 173.500 116.600 173.800 116.900 ;
        RECT 175.000 119.600 177.000 119.900 ;
        RECT 175.000 116.900 175.400 119.600 ;
        RECT 175.800 116.900 176.200 119.300 ;
        RECT 176.600 117.000 177.000 119.600 ;
        RECT 177.500 119.600 179.300 119.900 ;
        RECT 177.500 119.500 177.800 119.600 ;
        RECT 175.000 116.600 175.300 116.900 ;
        RECT 173.500 116.300 175.300 116.600 ;
        RECT 175.900 116.700 176.200 116.900 ;
        RECT 177.400 116.700 177.800 119.500 ;
        RECT 179.000 119.500 179.300 119.600 ;
        RECT 175.900 116.500 177.800 116.700 ;
        RECT 178.200 116.500 178.600 119.300 ;
        RECT 179.000 116.500 179.400 119.500 ;
        RECT 175.900 116.400 177.700 116.500 ;
        RECT 178.200 116.200 178.500 116.500 ;
        RECT 171.500 115.900 172.000 116.200 ;
        RECT 172.300 115.900 173.000 116.200 ;
        RECT 178.200 116.100 178.600 116.200 ;
        RECT 171.000 114.400 171.400 115.200 ;
        RECT 171.700 114.200 172.000 115.900 ;
        RECT 172.600 115.800 173.000 115.900 ;
        RECT 176.900 115.800 178.600 116.100 ;
        RECT 173.400 115.100 173.800 115.200 ;
        RECT 175.800 115.100 176.600 115.200 ;
        RECT 173.400 114.800 176.600 115.100 ;
        RECT 170.200 114.100 170.600 114.200 ;
        RECT 171.700 114.100 173.000 114.200 ;
        RECT 175.000 114.100 175.800 114.200 ;
        RECT 170.200 113.800 171.000 114.100 ;
        RECT 171.700 113.800 175.800 114.100 ;
        RECT 170.600 113.600 171.000 113.800 ;
        RECT 170.300 113.100 172.100 113.300 ;
        RECT 172.600 113.100 172.900 113.800 ;
        RECT 168.600 112.800 169.500 113.100 ;
        RECT 169.100 112.200 169.500 112.800 ;
        RECT 168.600 111.800 169.500 112.200 ;
        RECT 169.100 111.100 169.500 111.800 ;
        RECT 170.200 113.000 172.200 113.100 ;
        RECT 170.200 111.100 170.600 113.000 ;
        RECT 171.800 111.100 172.200 113.000 ;
        RECT 172.600 111.100 173.000 113.100 ;
        RECT 174.200 112.800 175.100 113.200 ;
        RECT 176.900 112.500 177.200 115.800 ;
        RECT 175.200 112.200 177.200 112.500 ;
        RECT 175.000 111.800 175.500 112.200 ;
        RECT 176.600 112.100 177.200 112.200 ;
        RECT 175.000 111.100 175.400 111.800 ;
        RECT 176.600 111.100 177.000 112.100 ;
        RECT 0.600 107.500 1.000 109.900 ;
        RECT 2.800 109.200 3.200 109.900 ;
        RECT 2.200 108.900 3.200 109.200 ;
        RECT 5.000 108.900 5.400 109.900 ;
        RECT 7.100 109.200 7.700 109.900 ;
        RECT 7.000 108.900 7.700 109.200 ;
        RECT 2.200 108.500 2.600 108.900 ;
        RECT 5.000 108.600 5.300 108.900 ;
        RECT 3.000 108.200 3.400 108.600 ;
        RECT 3.900 108.300 5.300 108.600 ;
        RECT 7.000 108.500 7.400 108.900 ;
        RECT 3.900 108.200 4.300 108.300 ;
        RECT 1.000 107.100 1.800 107.200 ;
        RECT 3.100 107.100 3.400 108.200 ;
        RECT 7.900 107.700 8.300 107.800 ;
        RECT 9.400 107.700 9.800 109.900 ;
        RECT 7.900 107.400 9.800 107.700 ;
        RECT 5.900 107.100 6.300 107.200 ;
        RECT 1.000 106.800 6.500 107.100 ;
        RECT 2.500 106.700 2.900 106.800 ;
        RECT 1.700 106.200 2.100 106.300 ;
        RECT 6.200 106.200 6.500 106.800 ;
        RECT 7.000 106.400 7.400 106.500 ;
        RECT 1.700 105.900 4.200 106.200 ;
        RECT 3.800 105.800 4.200 105.900 ;
        RECT 6.200 105.800 6.600 106.200 ;
        RECT 7.000 106.100 8.900 106.400 ;
        RECT 8.500 106.000 8.900 106.100 ;
        RECT 0.600 105.500 3.400 105.600 ;
        RECT 0.600 105.400 3.500 105.500 ;
        RECT 0.600 105.300 5.500 105.400 ;
        RECT 0.600 101.100 1.000 105.300 ;
        RECT 3.100 105.100 5.500 105.300 ;
        RECT 2.200 104.500 4.900 104.800 ;
        RECT 2.200 104.400 2.600 104.500 ;
        RECT 4.500 104.400 4.900 104.500 ;
        RECT 5.200 104.500 5.500 105.100 ;
        RECT 6.200 105.200 6.500 105.800 ;
        RECT 7.700 105.700 8.100 105.800 ;
        RECT 9.400 105.700 9.800 107.400 ;
        RECT 11.800 107.900 12.200 109.900 ;
        RECT 14.200 108.900 14.600 109.900 ;
        RECT 12.500 108.200 12.900 108.600 ;
        RECT 12.600 108.100 13.000 108.200 ;
        RECT 14.200 108.100 14.500 108.900 ;
        RECT 11.000 106.400 11.400 107.200 ;
        RECT 11.800 106.200 12.100 107.900 ;
        RECT 12.600 107.800 14.500 108.100 ;
        RECT 15.000 107.800 15.400 108.600 ;
        RECT 14.200 107.200 14.500 107.800 ;
        RECT 15.800 107.500 16.200 109.900 ;
        RECT 18.000 109.200 18.400 109.900 ;
        RECT 17.400 108.900 18.400 109.200 ;
        RECT 20.200 108.900 20.600 109.900 ;
        RECT 22.300 109.200 22.900 109.900 ;
        RECT 22.200 108.900 22.900 109.200 ;
        RECT 17.400 108.500 17.800 108.900 ;
        RECT 20.200 108.600 20.500 108.900 ;
        RECT 18.200 108.200 18.600 108.600 ;
        RECT 19.100 108.300 20.500 108.600 ;
        RECT 22.200 108.500 22.600 108.900 ;
        RECT 19.100 108.200 19.500 108.300 ;
        RECT 14.200 106.800 14.600 107.200 ;
        RECT 16.200 107.100 17.000 107.200 ;
        RECT 18.300 107.100 18.600 108.200 ;
        RECT 21.400 108.100 21.800 108.200 ;
        RECT 21.400 107.800 23.400 108.100 ;
        RECT 23.000 107.700 23.500 107.800 ;
        RECT 24.600 107.700 25.000 109.900 ;
        RECT 26.900 107.900 27.700 109.900 ;
        RECT 23.000 107.400 25.000 107.700 ;
        RECT 21.100 107.100 21.500 107.200 ;
        RECT 16.200 106.800 21.700 107.100 ;
        RECT 10.200 106.100 10.600 106.200 ;
        RECT 11.800 106.100 12.200 106.200 ;
        RECT 12.600 106.100 13.000 106.200 ;
        RECT 10.200 105.800 11.000 106.100 ;
        RECT 11.800 105.800 13.000 106.100 ;
        RECT 7.700 105.400 9.800 105.700 ;
        RECT 10.600 105.600 11.000 105.800 ;
        RECT 6.200 104.900 7.400 105.200 ;
        RECT 5.900 104.500 6.300 104.600 ;
        RECT 5.200 104.200 6.300 104.500 ;
        RECT 7.100 104.400 7.400 104.900 ;
        RECT 7.100 104.000 7.800 104.400 ;
        RECT 3.900 103.700 4.300 103.800 ;
        RECT 5.300 103.700 5.700 103.800 ;
        RECT 2.200 103.100 2.600 103.500 ;
        RECT 3.900 103.400 5.700 103.700 ;
        RECT 5.000 103.100 5.300 103.400 ;
        RECT 7.000 103.100 7.400 103.500 ;
        RECT 2.200 102.800 3.200 103.100 ;
        RECT 2.800 101.100 3.200 102.800 ;
        RECT 5.000 101.100 5.400 103.100 ;
        RECT 7.100 101.100 7.700 103.100 ;
        RECT 9.400 101.100 9.800 105.400 ;
        RECT 12.600 105.100 12.900 105.800 ;
        RECT 13.400 105.400 13.800 106.200 ;
        RECT 14.200 105.100 14.500 106.800 ;
        RECT 17.700 106.700 18.100 106.800 ;
        RECT 16.900 106.200 17.300 106.300 ;
        RECT 18.200 106.200 18.600 106.300 ;
        RECT 16.900 105.900 19.400 106.200 ;
        RECT 19.000 105.800 19.400 105.900 ;
        RECT 15.800 105.500 18.600 105.600 ;
        RECT 15.800 105.400 18.700 105.500 ;
        RECT 15.800 105.300 20.700 105.400 ;
        RECT 10.200 104.800 12.200 105.100 ;
        RECT 10.200 101.100 10.600 104.800 ;
        RECT 11.800 101.100 12.200 104.800 ;
        RECT 12.600 101.100 13.000 105.100 ;
        RECT 13.700 104.700 14.600 105.100 ;
        RECT 13.700 101.100 14.100 104.700 ;
        RECT 15.800 101.100 16.200 105.300 ;
        RECT 18.300 105.100 20.700 105.300 ;
        RECT 17.400 104.500 20.100 104.800 ;
        RECT 17.400 104.400 17.800 104.500 ;
        RECT 19.700 104.400 20.100 104.500 ;
        RECT 20.400 104.500 20.700 105.100 ;
        RECT 21.400 105.200 21.700 106.800 ;
        RECT 22.200 106.400 22.600 106.500 ;
        RECT 22.200 106.100 24.100 106.400 ;
        RECT 23.700 106.000 24.100 106.100 ;
        RECT 24.600 106.100 25.000 107.400 ;
        RECT 26.200 106.400 26.600 107.200 ;
        RECT 27.100 106.200 27.400 107.900 ;
        RECT 29.400 107.500 29.800 109.900 ;
        RECT 31.600 109.200 32.000 109.900 ;
        RECT 31.000 108.900 32.000 109.200 ;
        RECT 33.800 108.900 34.200 109.900 ;
        RECT 35.900 109.200 36.500 109.900 ;
        RECT 35.800 108.900 36.500 109.200 ;
        RECT 31.000 108.500 31.400 108.900 ;
        RECT 33.800 108.600 34.100 108.900 ;
        RECT 31.800 108.200 32.200 108.600 ;
        RECT 32.700 108.300 34.100 108.600 ;
        RECT 35.800 108.500 36.200 108.900 ;
        RECT 32.700 108.200 33.100 108.300 ;
        RECT 27.800 106.800 28.200 107.200 ;
        RECT 29.800 107.100 30.600 107.200 ;
        RECT 31.900 107.100 32.200 108.200 ;
        RECT 36.700 107.700 37.100 107.800 ;
        RECT 38.200 107.700 38.600 109.900 ;
        RECT 36.700 107.400 38.600 107.700 ;
        RECT 34.700 107.100 35.100 107.200 ;
        RECT 29.800 106.800 35.300 107.100 ;
        RECT 27.800 106.600 28.100 106.800 ;
        RECT 31.300 106.700 31.700 106.800 ;
        RECT 27.700 106.200 28.100 106.600 ;
        RECT 30.500 106.200 30.900 106.300 ;
        RECT 25.400 106.100 25.800 106.200 ;
        RECT 24.600 105.800 26.200 106.100 ;
        RECT 27.000 105.800 27.400 106.200 ;
        RECT 22.900 105.700 23.300 105.800 ;
        RECT 24.600 105.700 25.000 105.800 ;
        RECT 22.900 105.400 25.000 105.700 ;
        RECT 25.800 105.600 26.200 105.800 ;
        RECT 27.100 105.700 27.400 105.800 ;
        RECT 27.100 105.400 28.100 105.700 ;
        RECT 28.600 105.400 29.000 106.200 ;
        RECT 30.500 105.900 33.000 106.200 ;
        RECT 32.600 105.800 33.000 105.900 ;
        RECT 29.400 105.500 32.200 105.600 ;
        RECT 29.400 105.400 32.300 105.500 ;
        RECT 21.400 104.900 22.600 105.200 ;
        RECT 21.100 104.500 21.500 104.600 ;
        RECT 20.400 104.200 21.500 104.500 ;
        RECT 22.300 104.400 22.600 104.900 ;
        RECT 22.300 104.000 23.000 104.400 ;
        RECT 19.100 103.700 19.500 103.800 ;
        RECT 20.500 103.700 20.900 103.800 ;
        RECT 17.400 103.100 17.800 103.500 ;
        RECT 19.100 103.400 20.900 103.700 ;
        RECT 20.200 103.100 20.500 103.400 ;
        RECT 22.200 103.100 22.600 103.500 ;
        RECT 17.400 102.800 18.400 103.100 ;
        RECT 18.000 101.100 18.400 102.800 ;
        RECT 20.200 101.100 20.600 103.100 ;
        RECT 22.300 101.100 22.900 103.100 ;
        RECT 24.600 101.100 25.000 105.400 ;
        RECT 27.800 105.100 28.100 105.400 ;
        RECT 29.400 105.300 34.300 105.400 ;
        RECT 25.400 104.800 27.400 105.100 ;
        RECT 25.400 101.100 25.800 104.800 ;
        RECT 27.000 101.400 27.400 104.800 ;
        RECT 27.800 101.700 28.200 105.100 ;
        RECT 28.600 101.400 29.000 105.100 ;
        RECT 27.000 101.100 29.000 101.400 ;
        RECT 29.400 101.100 29.800 105.300 ;
        RECT 31.900 105.100 34.300 105.300 ;
        RECT 31.000 104.500 33.700 104.800 ;
        RECT 31.000 104.400 31.400 104.500 ;
        RECT 33.300 104.400 33.700 104.500 ;
        RECT 34.000 104.500 34.300 105.100 ;
        RECT 35.000 105.200 35.300 106.800 ;
        RECT 35.800 106.400 36.200 106.500 ;
        RECT 35.800 106.100 37.700 106.400 ;
        RECT 37.300 106.000 37.700 106.100 ;
        RECT 36.500 105.700 36.900 105.800 ;
        RECT 38.200 105.700 38.600 107.400 ;
        RECT 40.600 108.500 41.000 109.500 ;
        RECT 40.600 107.400 40.900 108.500 ;
        RECT 42.700 108.000 43.100 109.500 ;
        RECT 42.700 107.700 43.500 108.000 ;
        RECT 43.100 107.500 43.500 107.700 ;
        RECT 40.600 107.100 42.700 107.400 ;
        RECT 42.200 106.900 42.700 107.100 ;
        RECT 43.200 107.200 43.500 107.500 ;
        RECT 39.800 106.100 40.200 106.200 ;
        RECT 40.600 106.100 41.000 106.600 ;
        RECT 39.800 105.800 41.000 106.100 ;
        RECT 41.400 105.800 41.800 106.600 ;
        RECT 42.200 106.500 42.900 106.900 ;
        RECT 43.200 106.800 44.200 107.200 ;
        RECT 36.500 105.400 38.600 105.700 ;
        RECT 42.200 105.500 42.500 106.500 ;
        RECT 35.000 104.900 36.200 105.200 ;
        RECT 34.700 104.500 35.100 104.600 ;
        RECT 34.000 104.200 35.100 104.500 ;
        RECT 35.900 104.400 36.200 104.900 ;
        RECT 35.900 104.000 36.600 104.400 ;
        RECT 32.700 103.700 33.100 103.800 ;
        RECT 34.100 103.700 34.500 103.800 ;
        RECT 31.000 103.100 31.400 103.500 ;
        RECT 32.700 103.400 34.500 103.700 ;
        RECT 33.800 103.100 34.100 103.400 ;
        RECT 35.800 103.100 36.200 103.500 ;
        RECT 31.000 102.800 32.000 103.100 ;
        RECT 31.600 101.100 32.000 102.800 ;
        RECT 33.800 101.100 34.200 103.100 ;
        RECT 35.900 101.100 36.500 103.100 ;
        RECT 38.200 101.100 38.600 105.400 ;
        RECT 40.600 105.200 42.500 105.500 ;
        RECT 43.200 105.200 43.500 106.800 ;
        RECT 43.800 106.100 44.200 106.200 ;
        RECT 45.400 106.100 45.800 109.900 ;
        RECT 46.200 107.800 46.600 108.600 ;
        RECT 48.300 108.200 48.700 109.900 ;
        RECT 47.800 107.900 48.700 108.200 ;
        RECT 50.000 109.100 50.400 109.900 ;
        RECT 51.000 109.100 51.400 109.200 ;
        RECT 50.000 108.800 51.400 109.100 ;
        RECT 47.000 106.800 47.400 107.600 ;
        RECT 43.800 105.800 45.800 106.100 ;
        RECT 43.800 105.400 44.200 105.800 ;
        RECT 40.600 103.500 40.900 105.200 ;
        RECT 43.000 104.900 43.500 105.200 ;
        RECT 42.700 104.600 43.500 104.900 ;
        RECT 40.600 101.500 41.000 103.500 ;
        RECT 42.700 101.100 43.100 104.600 ;
        RECT 45.400 101.100 45.800 105.800 ;
        RECT 47.000 105.100 47.400 105.200 ;
        RECT 47.800 105.100 48.200 107.900 ;
        RECT 50.000 107.100 50.400 108.800 ;
        RECT 53.900 107.900 54.700 109.900 ;
        RECT 57.400 108.900 57.800 109.900 ;
        RECT 49.500 106.900 50.400 107.100 ;
        RECT 49.500 106.800 50.300 106.900 ;
        RECT 53.400 106.800 53.800 107.200 ;
        RECT 49.500 105.200 49.800 106.800 ;
        RECT 53.500 106.600 53.800 106.800 ;
        RECT 53.500 106.200 53.900 106.600 ;
        RECT 54.200 106.200 54.500 107.900 ;
        RECT 57.400 107.200 57.700 108.900 ;
        RECT 58.200 107.800 58.600 108.600 ;
        RECT 59.100 108.200 59.500 108.600 ;
        RECT 59.000 107.800 59.400 108.200 ;
        RECT 59.800 107.900 60.200 109.900 ;
        RECT 55.000 106.400 55.400 107.200 ;
        RECT 57.400 107.100 57.800 107.200 ;
        RECT 59.000 107.100 59.300 107.800 ;
        RECT 57.400 106.800 59.300 107.100 ;
        RECT 50.200 105.800 51.400 106.200 ;
        RECT 47.000 104.800 48.200 105.100 ;
        RECT 47.800 101.100 48.200 104.800 ;
        RECT 48.600 104.400 49.000 105.200 ;
        RECT 49.400 104.800 49.800 105.200 ;
        RECT 51.800 104.800 52.200 105.600 ;
        RECT 52.600 105.400 53.000 106.200 ;
        RECT 54.200 105.800 54.600 106.200 ;
        RECT 55.800 106.100 56.200 106.200 ;
        RECT 55.400 105.800 56.200 106.100 ;
        RECT 54.200 105.700 54.500 105.800 ;
        RECT 53.500 105.400 54.500 105.700 ;
        RECT 55.400 105.600 55.800 105.800 ;
        RECT 56.600 105.400 57.000 106.200 ;
        RECT 53.500 105.100 53.800 105.400 ;
        RECT 57.400 105.100 57.700 106.800 ;
        RECT 59.000 106.100 59.400 106.200 ;
        RECT 59.900 106.100 60.200 107.900 ;
        RECT 60.600 106.400 61.000 107.200 ;
        RECT 64.000 107.100 64.400 109.900 ;
        RECT 65.700 108.200 66.100 109.900 ;
        RECT 65.700 107.900 66.600 108.200 ;
        RECT 64.000 106.900 64.900 107.100 ;
        RECT 64.100 106.800 64.900 106.900 ;
        RECT 61.400 106.100 61.800 106.200 ;
        RECT 59.000 105.800 60.200 106.100 ;
        RECT 61.000 105.800 61.800 106.100 ;
        RECT 63.000 105.800 63.800 106.200 ;
        RECT 59.100 105.100 59.400 105.800 ;
        RECT 61.000 105.600 61.400 105.800 ;
        RECT 49.500 103.500 49.800 104.800 ;
        RECT 50.200 103.800 50.600 104.600 ;
        RECT 49.500 103.200 51.300 103.500 ;
        RECT 49.500 103.100 49.800 103.200 ;
        RECT 49.400 101.100 49.800 103.100 ;
        RECT 51.000 103.100 51.300 103.200 ;
        RECT 51.000 101.100 51.400 103.100 ;
        RECT 52.600 101.400 53.000 105.100 ;
        RECT 53.400 101.700 53.800 105.100 ;
        RECT 54.200 104.800 56.200 105.100 ;
        RECT 54.200 101.400 54.600 104.800 ;
        RECT 52.600 101.100 54.600 101.400 ;
        RECT 55.800 101.100 56.200 104.800 ;
        RECT 56.900 104.700 57.800 105.100 ;
        RECT 56.900 101.100 57.300 104.700 ;
        RECT 59.000 101.100 59.400 105.100 ;
        RECT 59.800 104.800 61.800 105.100 ;
        RECT 62.200 104.800 62.600 105.600 ;
        RECT 64.600 105.200 64.900 106.800 ;
        RECT 65.400 106.800 65.800 107.200 ;
        RECT 65.400 106.100 65.700 106.800 ;
        RECT 66.200 106.100 66.600 107.900 ;
        RECT 67.800 107.700 68.200 109.900 ;
        RECT 69.900 109.200 70.500 109.900 ;
        RECT 69.900 108.900 70.600 109.200 ;
        RECT 72.200 108.900 72.600 109.900 ;
        RECT 74.400 109.200 74.800 109.900 ;
        RECT 74.400 108.900 75.400 109.200 ;
        RECT 70.200 108.500 70.600 108.900 ;
        RECT 72.300 108.600 72.600 108.900 ;
        RECT 72.300 108.300 73.700 108.600 ;
        RECT 73.300 108.200 73.700 108.300 ;
        RECT 74.200 108.200 74.600 108.600 ;
        RECT 75.000 108.500 75.400 108.900 ;
        RECT 69.300 107.700 69.700 107.800 ;
        RECT 67.000 106.800 67.400 107.600 ;
        RECT 67.800 107.400 69.700 107.700 ;
        RECT 65.400 105.800 66.600 106.100 ;
        RECT 64.600 104.800 65.000 105.200 ;
        RECT 59.800 101.100 60.200 104.800 ;
        RECT 61.400 101.100 61.800 104.800 ;
        RECT 63.800 103.800 64.200 104.600 ;
        RECT 64.600 103.500 64.900 104.800 ;
        RECT 65.400 104.400 65.800 105.200 ;
        RECT 63.100 103.200 64.900 103.500 ;
        RECT 63.100 103.100 63.400 103.200 ;
        RECT 63.000 101.100 63.400 103.100 ;
        RECT 64.600 103.100 64.900 103.200 ;
        RECT 64.600 101.100 65.000 103.100 ;
        RECT 66.200 101.100 66.600 105.800 ;
        RECT 67.800 105.700 68.200 107.400 ;
        RECT 71.300 107.100 71.700 107.200 ;
        RECT 74.200 107.100 74.500 108.200 ;
        RECT 76.600 107.500 77.000 109.900 ;
        RECT 79.000 109.200 79.400 109.900 ;
        RECT 79.000 108.900 79.500 109.200 ;
        RECT 79.200 108.800 79.500 108.900 ;
        RECT 80.600 108.900 81.000 109.900 ;
        RECT 80.600 108.800 81.200 108.900 ;
        RECT 79.200 108.500 81.200 108.800 ;
        RECT 78.200 107.800 79.100 108.200 ;
        RECT 75.800 107.100 76.600 107.200 ;
        RECT 71.100 106.800 76.600 107.100 ;
        RECT 78.200 107.100 78.600 107.200 ;
        RECT 79.000 107.100 79.800 107.200 ;
        RECT 78.200 106.800 79.800 107.100 ;
        RECT 80.900 107.100 81.200 108.500 ;
        RECT 82.200 107.800 82.600 108.200 ;
        RECT 85.300 107.900 86.100 109.900 ;
        RECT 88.100 109.200 88.500 109.900 ;
        RECT 87.800 108.800 88.500 109.200 ;
        RECT 88.100 108.200 88.500 108.800 ;
        RECT 88.100 107.900 89.000 108.200 ;
        RECT 82.200 107.100 82.500 107.800 ;
        RECT 80.900 106.800 82.500 107.100 ;
        RECT 83.000 107.100 83.400 107.200 ;
        RECT 84.600 107.100 85.000 107.200 ;
        RECT 83.000 106.800 85.000 107.100 ;
        RECT 70.200 106.400 70.600 106.500 ;
        RECT 68.700 106.100 70.600 106.400 ;
        RECT 68.700 106.000 69.100 106.100 ;
        RECT 69.500 105.700 69.900 105.800 ;
        RECT 67.800 105.400 69.900 105.700 ;
        RECT 67.800 101.100 68.200 105.400 ;
        RECT 71.100 105.200 71.400 106.800 ;
        RECT 74.700 106.700 75.100 106.800 ;
        RECT 75.500 106.200 75.900 106.300 ;
        RECT 71.800 106.100 72.200 106.200 ;
        RECT 73.400 106.100 75.900 106.200 ;
        RECT 71.800 105.900 75.900 106.100 ;
        RECT 71.800 105.800 73.800 105.900 ;
        RECT 79.800 105.800 80.600 106.200 ;
        RECT 74.200 105.500 77.000 105.600 ;
        RECT 74.100 105.400 77.000 105.500 ;
        RECT 70.200 104.900 71.400 105.200 ;
        RECT 72.100 105.300 77.000 105.400 ;
        RECT 72.100 105.100 74.500 105.300 ;
        RECT 70.200 104.400 70.500 104.900 ;
        RECT 69.800 104.200 70.500 104.400 ;
        RECT 71.300 104.500 71.700 104.600 ;
        RECT 72.100 104.500 72.400 105.100 ;
        RECT 71.300 104.200 72.400 104.500 ;
        RECT 72.700 104.500 75.400 104.800 ;
        RECT 72.700 104.400 73.100 104.500 ;
        RECT 75.000 104.400 75.400 104.500 ;
        RECT 69.400 104.000 70.500 104.200 ;
        RECT 69.400 103.800 70.100 104.000 ;
        RECT 71.900 103.700 72.300 103.800 ;
        RECT 73.300 103.700 73.700 103.800 ;
        RECT 70.200 103.100 70.600 103.500 ;
        RECT 71.900 103.400 73.700 103.700 ;
        RECT 72.300 103.100 72.600 103.400 ;
        RECT 75.000 103.100 75.400 103.500 ;
        RECT 69.900 101.100 70.500 103.100 ;
        RECT 72.200 101.100 72.600 103.100 ;
        RECT 74.400 102.800 75.400 103.100 ;
        RECT 74.400 101.100 74.800 102.800 ;
        RECT 76.600 101.100 77.000 105.300 ;
        RECT 80.900 105.200 81.200 106.800 ;
        RECT 84.600 106.400 85.000 106.800 ;
        RECT 85.500 106.200 85.800 107.900 ;
        RECT 86.200 106.800 86.600 107.200 ;
        RECT 86.200 106.600 86.500 106.800 ;
        RECT 86.100 106.200 86.500 106.600 ;
        RECT 82.200 106.100 82.600 106.200 ;
        RECT 83.800 106.100 84.200 106.200 ;
        RECT 82.200 105.800 84.600 106.100 ;
        RECT 85.400 105.800 85.800 106.200 ;
        RECT 84.200 105.600 84.600 105.800 ;
        RECT 85.500 105.700 85.800 105.800 ;
        RECT 85.500 105.400 86.500 105.700 ;
        RECT 87.000 105.400 87.400 106.200 ;
        RECT 80.900 104.900 82.600 105.200 ;
        RECT 86.200 105.100 86.500 105.400 ;
        RECT 82.200 104.800 82.600 104.900 ;
        RECT 83.800 104.800 85.800 105.100 ;
        RECT 77.500 104.400 79.300 104.700 ;
        RECT 77.500 104.100 77.800 104.400 ;
        RECT 77.400 101.100 77.800 104.100 ;
        RECT 79.000 104.100 79.300 104.400 ;
        RECT 79.900 104.500 81.700 104.600 ;
        RECT 82.200 104.500 82.500 104.800 ;
        RECT 79.900 104.300 81.800 104.500 ;
        RECT 79.900 104.100 80.200 104.300 ;
        RECT 79.000 101.400 79.400 104.100 ;
        RECT 79.800 101.700 80.200 104.100 ;
        RECT 80.600 101.400 81.000 104.000 ;
        RECT 81.400 101.500 81.800 104.300 ;
        RECT 82.200 101.700 82.600 104.500 ;
        RECT 79.000 101.100 81.000 101.400 ;
        RECT 81.500 101.400 81.800 101.500 ;
        RECT 83.000 101.500 83.400 104.500 ;
        RECT 83.000 101.400 83.300 101.500 ;
        RECT 81.500 101.100 83.300 101.400 ;
        RECT 83.800 101.100 84.200 104.800 ;
        RECT 85.400 101.400 85.800 104.800 ;
        RECT 86.200 101.700 86.600 105.100 ;
        RECT 87.000 101.400 87.400 105.100 ;
        RECT 87.800 104.400 88.200 105.200 ;
        RECT 85.400 101.100 87.400 101.400 ;
        RECT 88.600 101.100 89.000 107.900 ;
        RECT 92.600 107.600 93.000 109.900 ;
        RECT 94.200 107.600 94.600 109.900 ;
        RECT 95.800 107.600 96.200 109.900 ;
        RECT 97.400 107.600 97.800 109.900 ;
        RECT 100.500 107.900 101.300 109.900 ;
        RECT 89.400 107.100 89.800 107.600 ;
        RECT 91.800 107.200 93.000 107.600 ;
        RECT 93.500 107.200 94.600 107.600 ;
        RECT 95.100 107.200 96.200 107.600 ;
        RECT 96.900 107.200 97.800 107.600 ;
        RECT 91.000 107.100 91.400 107.200 ;
        RECT 89.400 106.800 91.400 107.100 ;
        RECT 91.800 105.800 92.200 107.200 ;
        RECT 93.500 106.900 93.900 107.200 ;
        RECT 95.100 106.900 95.500 107.200 ;
        RECT 96.900 106.900 97.300 107.200 ;
        RECT 92.600 106.500 93.900 106.900 ;
        RECT 94.300 106.500 95.500 106.900 ;
        RECT 96.000 106.500 97.300 106.900 ;
        RECT 93.500 105.800 93.900 106.500 ;
        RECT 95.100 105.800 95.500 106.500 ;
        RECT 96.900 105.800 97.300 106.500 ;
        RECT 99.800 106.400 100.200 107.200 ;
        RECT 100.700 106.200 101.000 107.900 ;
        RECT 101.400 106.800 101.800 107.200 ;
        RECT 103.000 106.800 103.400 107.600 ;
        RECT 101.400 106.600 101.700 106.800 ;
        RECT 101.300 106.200 101.700 106.600 ;
        RECT 99.000 106.100 99.400 106.200 ;
        RECT 99.000 105.800 99.800 106.100 ;
        RECT 100.600 105.800 101.000 106.200 ;
        RECT 91.800 105.400 93.000 105.800 ;
        RECT 93.500 105.400 94.600 105.800 ;
        RECT 95.100 105.400 96.200 105.800 ;
        RECT 96.900 105.400 97.800 105.800 ;
        RECT 99.400 105.600 99.800 105.800 ;
        RECT 100.700 105.700 101.000 105.800 ;
        RECT 100.700 105.400 101.700 105.700 ;
        RECT 102.200 105.400 102.600 106.200 ;
        RECT 92.600 101.100 93.000 105.400 ;
        RECT 94.200 101.100 94.600 105.400 ;
        RECT 95.800 101.100 96.200 105.400 ;
        RECT 97.400 101.100 97.800 105.400 ;
        RECT 101.400 105.100 101.700 105.400 ;
        RECT 99.000 104.800 101.000 105.100 ;
        RECT 99.000 101.100 99.400 104.800 ;
        RECT 100.600 101.400 101.000 104.800 ;
        RECT 101.400 101.700 101.800 105.100 ;
        RECT 102.200 101.400 102.600 105.100 ;
        RECT 100.600 101.100 102.600 101.400 ;
        RECT 103.800 101.100 104.200 109.900 ;
        RECT 106.900 107.900 107.700 109.900 ;
        RECT 106.200 106.400 106.600 107.200 ;
        RECT 107.100 106.200 107.400 107.900 ;
        RECT 109.400 107.800 109.800 108.600 ;
        RECT 107.800 106.800 108.200 107.200 ;
        RECT 107.800 106.600 108.100 106.800 ;
        RECT 107.700 106.200 108.100 106.600 ;
        RECT 104.600 106.100 105.000 106.200 ;
        RECT 105.400 106.100 105.800 106.200 ;
        RECT 104.600 105.800 106.200 106.100 ;
        RECT 107.000 105.800 107.400 106.200 ;
        RECT 105.800 105.600 106.200 105.800 ;
        RECT 107.100 105.700 107.400 105.800 ;
        RECT 108.600 106.100 109.000 106.200 ;
        RECT 109.400 106.100 109.800 106.200 ;
        RECT 108.600 105.800 109.800 106.100 ;
        RECT 107.100 105.400 108.100 105.700 ;
        RECT 108.600 105.400 109.000 105.800 ;
        RECT 107.800 105.100 108.100 105.400 ;
        RECT 105.400 104.800 107.400 105.100 ;
        RECT 105.400 101.100 105.800 104.800 ;
        RECT 107.000 101.400 107.400 104.800 ;
        RECT 107.800 101.700 108.200 105.100 ;
        RECT 108.600 101.400 109.000 105.100 ;
        RECT 107.000 101.100 109.000 101.400 ;
        RECT 110.200 101.100 110.600 109.900 ;
        RECT 111.000 107.700 111.400 109.900 ;
        RECT 113.100 109.200 113.700 109.900 ;
        RECT 113.100 108.900 113.800 109.200 ;
        RECT 115.400 108.900 115.800 109.900 ;
        RECT 117.600 109.200 118.000 109.900 ;
        RECT 117.600 108.900 118.600 109.200 ;
        RECT 113.400 108.500 113.800 108.900 ;
        RECT 115.500 108.600 115.800 108.900 ;
        RECT 115.500 108.300 116.900 108.600 ;
        RECT 116.500 108.200 116.900 108.300 ;
        RECT 117.400 108.200 117.800 108.600 ;
        RECT 118.200 108.500 118.600 108.900 ;
        RECT 112.500 107.700 112.900 107.800 ;
        RECT 111.000 107.400 112.900 107.700 ;
        RECT 111.000 105.700 111.400 107.400 ;
        RECT 114.500 107.100 114.900 107.200 ;
        RECT 117.400 107.100 117.700 108.200 ;
        RECT 119.800 107.500 120.200 109.900 ;
        RECT 120.600 107.500 121.000 109.900 ;
        RECT 122.800 109.200 123.200 109.900 ;
        RECT 122.200 108.900 123.200 109.200 ;
        RECT 125.000 108.900 125.400 109.900 ;
        RECT 127.100 109.200 127.700 109.900 ;
        RECT 127.000 108.900 127.700 109.200 ;
        RECT 122.200 108.500 122.600 108.900 ;
        RECT 125.000 108.600 125.300 108.900 ;
        RECT 123.000 108.200 123.400 108.600 ;
        RECT 123.900 108.300 125.300 108.600 ;
        RECT 127.000 108.500 127.400 108.900 ;
        RECT 123.900 108.200 124.300 108.300 ;
        RECT 119.000 107.100 119.800 107.200 ;
        RECT 121.000 107.100 121.800 107.200 ;
        RECT 123.100 107.100 123.400 108.200 ;
        RECT 127.900 107.700 128.300 107.800 ;
        RECT 129.400 107.700 129.800 109.900 ;
        RECT 127.900 107.400 129.800 107.700 ;
        RECT 130.200 107.500 130.600 109.900 ;
        RECT 132.400 109.200 132.800 109.900 ;
        RECT 131.800 108.900 132.800 109.200 ;
        RECT 134.600 108.900 135.000 109.900 ;
        RECT 136.700 109.200 137.300 109.900 ;
        RECT 136.600 108.900 137.300 109.200 ;
        RECT 139.000 109.100 139.400 109.900 ;
        RECT 131.800 108.500 132.200 108.900 ;
        RECT 134.600 108.600 134.900 108.900 ;
        RECT 132.600 108.200 133.000 108.600 ;
        RECT 133.500 108.300 134.900 108.600 ;
        RECT 136.600 108.500 137.000 108.900 ;
        RECT 139.000 108.800 140.100 109.100 ;
        RECT 133.500 108.200 133.900 108.300 ;
        RECT 125.900 107.100 126.300 107.200 ;
        RECT 114.300 106.800 126.500 107.100 ;
        RECT 113.400 106.400 113.800 106.500 ;
        RECT 111.900 106.100 113.800 106.400 ;
        RECT 111.900 106.000 112.300 106.100 ;
        RECT 112.700 105.700 113.100 105.800 ;
        RECT 111.000 105.400 113.100 105.700 ;
        RECT 111.000 101.100 111.400 105.400 ;
        RECT 114.300 105.200 114.600 106.800 ;
        RECT 117.900 106.700 118.300 106.800 ;
        RECT 122.500 106.700 122.900 106.800 ;
        RECT 118.700 106.200 119.100 106.300 ;
        RECT 116.600 105.900 119.100 106.200 ;
        RECT 121.700 106.200 122.100 106.300 ;
        RECT 123.000 106.200 123.400 106.300 ;
        RECT 126.200 106.200 126.500 106.800 ;
        RECT 127.000 106.400 127.400 106.500 ;
        RECT 121.700 105.900 124.200 106.200 ;
        RECT 116.600 105.800 117.000 105.900 ;
        RECT 123.800 105.800 124.200 105.900 ;
        RECT 126.200 105.800 126.600 106.200 ;
        RECT 127.000 106.100 128.900 106.400 ;
        RECT 128.500 106.000 128.900 106.100 ;
        RECT 117.400 105.500 120.200 105.600 ;
        RECT 117.300 105.400 120.200 105.500 ;
        RECT 113.400 104.900 114.600 105.200 ;
        RECT 115.300 105.300 120.200 105.400 ;
        RECT 115.300 105.100 117.700 105.300 ;
        RECT 113.400 104.400 113.700 104.900 ;
        RECT 113.000 104.000 113.700 104.400 ;
        RECT 114.500 104.500 114.900 104.600 ;
        RECT 115.300 104.500 115.600 105.100 ;
        RECT 114.500 104.200 115.600 104.500 ;
        RECT 115.900 104.500 118.600 104.800 ;
        RECT 115.900 104.400 116.300 104.500 ;
        RECT 118.200 104.400 118.600 104.500 ;
        RECT 115.100 103.700 115.500 103.800 ;
        RECT 116.500 103.700 116.900 103.800 ;
        RECT 113.400 103.100 113.800 103.500 ;
        RECT 115.100 103.400 116.900 103.700 ;
        RECT 115.500 103.100 115.800 103.400 ;
        RECT 118.200 103.100 118.600 103.500 ;
        RECT 113.100 101.100 113.700 103.100 ;
        RECT 115.400 101.100 115.800 103.100 ;
        RECT 117.600 102.800 118.600 103.100 ;
        RECT 117.600 101.100 118.000 102.800 ;
        RECT 119.800 101.100 120.200 105.300 ;
        RECT 120.600 105.500 123.400 105.600 ;
        RECT 120.600 105.400 123.500 105.500 ;
        RECT 120.600 105.300 125.500 105.400 ;
        RECT 120.600 101.100 121.000 105.300 ;
        RECT 123.100 105.100 125.500 105.300 ;
        RECT 122.200 104.500 124.900 104.800 ;
        RECT 122.200 104.400 122.600 104.500 ;
        RECT 124.500 104.400 124.900 104.500 ;
        RECT 125.200 104.500 125.500 105.100 ;
        RECT 126.200 105.200 126.500 105.800 ;
        RECT 127.700 105.700 128.100 105.800 ;
        RECT 129.400 105.700 129.800 107.400 ;
        RECT 130.600 107.100 131.400 107.200 ;
        RECT 132.700 107.100 133.000 108.200 ;
        RECT 137.500 107.700 137.900 107.800 ;
        RECT 139.000 107.700 139.400 108.800 ;
        RECT 139.800 108.100 140.100 108.800 ;
        RECT 141.400 108.100 141.800 108.600 ;
        RECT 139.800 107.800 141.800 108.100 ;
        RECT 137.500 107.400 139.400 107.700 ;
        RECT 135.500 107.100 136.200 107.200 ;
        RECT 130.600 106.800 136.200 107.100 ;
        RECT 132.100 106.700 132.500 106.800 ;
        RECT 131.300 106.200 131.700 106.300 ;
        RECT 131.300 106.100 133.800 106.200 ;
        RECT 134.200 106.100 134.600 106.200 ;
        RECT 131.300 105.900 134.600 106.100 ;
        RECT 133.400 105.800 134.600 105.900 ;
        RECT 127.700 105.400 129.800 105.700 ;
        RECT 126.200 104.900 127.400 105.200 ;
        RECT 125.900 104.500 126.300 104.600 ;
        RECT 125.200 104.200 126.300 104.500 ;
        RECT 127.100 104.400 127.400 104.900 ;
        RECT 127.100 104.000 127.800 104.400 ;
        RECT 123.900 103.700 124.300 103.800 ;
        RECT 125.300 103.700 125.700 103.800 ;
        RECT 122.200 103.100 122.600 103.500 ;
        RECT 123.900 103.400 125.700 103.700 ;
        RECT 125.000 103.100 125.300 103.400 ;
        RECT 127.000 103.100 127.400 103.500 ;
        RECT 122.200 102.800 123.200 103.100 ;
        RECT 122.800 101.100 123.200 102.800 ;
        RECT 125.000 101.100 125.400 103.100 ;
        RECT 127.100 101.100 127.700 103.100 ;
        RECT 129.400 101.100 129.800 105.400 ;
        RECT 130.200 105.500 133.000 105.600 ;
        RECT 130.200 105.400 133.100 105.500 ;
        RECT 130.200 105.300 135.100 105.400 ;
        RECT 130.200 101.100 130.600 105.300 ;
        RECT 132.700 105.100 135.100 105.300 ;
        RECT 131.800 104.500 134.500 104.800 ;
        RECT 131.800 104.400 132.200 104.500 ;
        RECT 134.100 104.400 134.500 104.500 ;
        RECT 134.800 104.500 135.100 105.100 ;
        RECT 135.800 105.200 136.100 106.800 ;
        RECT 136.600 106.400 137.000 106.500 ;
        RECT 136.600 106.100 138.500 106.400 ;
        RECT 138.100 106.000 138.500 106.100 ;
        RECT 137.300 105.700 137.700 105.800 ;
        RECT 139.000 105.700 139.400 107.400 ;
        RECT 137.300 105.400 139.400 105.700 ;
        RECT 135.800 104.900 137.000 105.200 ;
        RECT 135.500 104.500 135.900 104.600 ;
        RECT 134.800 104.200 135.900 104.500 ;
        RECT 136.700 104.400 137.000 104.900 ;
        RECT 136.700 104.000 137.400 104.400 ;
        RECT 133.500 103.700 133.900 103.800 ;
        RECT 134.900 103.700 135.300 103.800 ;
        RECT 131.800 103.100 132.200 103.500 ;
        RECT 133.500 103.400 135.300 103.700 ;
        RECT 134.600 103.100 134.900 103.400 ;
        RECT 136.600 103.100 137.000 103.500 ;
        RECT 131.800 102.800 132.800 103.100 ;
        RECT 132.400 101.100 132.800 102.800 ;
        RECT 134.600 101.100 135.000 103.100 ;
        RECT 136.700 101.100 137.300 103.100 ;
        RECT 139.000 101.100 139.400 105.400 ;
        RECT 142.200 107.100 142.600 109.900 ;
        RECT 144.900 108.000 145.300 109.500 ;
        RECT 147.000 108.500 147.400 109.500 ;
        RECT 144.500 107.700 145.300 108.000 ;
        RECT 144.500 107.500 144.900 107.700 ;
        RECT 144.500 107.200 144.800 107.500 ;
        RECT 147.100 107.400 147.400 108.500 ;
        RECT 147.800 107.800 148.200 108.600 ;
        RECT 142.200 106.800 143.300 107.100 ;
        RECT 143.800 106.800 144.800 107.200 ;
        RECT 145.300 107.100 147.400 107.400 ;
        RECT 145.300 106.900 145.800 107.100 ;
        RECT 142.200 101.100 142.600 106.800 ;
        RECT 143.000 106.200 143.300 106.800 ;
        RECT 143.000 105.800 143.400 106.200 ;
        RECT 143.800 105.400 144.200 106.200 ;
        RECT 144.500 104.900 144.800 106.800 ;
        RECT 145.100 106.500 145.800 106.900 ;
        RECT 145.500 105.500 145.800 106.500 ;
        RECT 146.200 105.800 146.600 106.600 ;
        RECT 147.000 105.800 147.400 106.600 ;
        RECT 147.800 106.100 148.200 106.200 ;
        RECT 148.600 106.100 149.000 109.900 ;
        RECT 147.800 105.800 149.000 106.100 ;
        RECT 145.500 105.200 147.400 105.500 ;
        RECT 144.500 104.600 145.300 104.900 ;
        RECT 144.900 101.100 145.300 104.600 ;
        RECT 147.100 103.500 147.400 105.200 ;
        RECT 147.000 101.500 147.400 103.500 ;
        RECT 148.600 101.100 149.000 105.800 ;
        RECT 149.400 107.700 149.800 109.900 ;
        RECT 151.500 109.200 152.100 109.900 ;
        RECT 151.500 108.900 152.200 109.200 ;
        RECT 153.800 108.900 154.200 109.900 ;
        RECT 156.000 109.200 156.400 109.900 ;
        RECT 156.000 108.900 157.000 109.200 ;
        RECT 151.800 108.500 152.200 108.900 ;
        RECT 153.900 108.600 154.200 108.900 ;
        RECT 153.900 108.300 155.300 108.600 ;
        RECT 154.900 108.200 155.300 108.300 ;
        RECT 155.800 107.800 156.200 108.600 ;
        RECT 156.600 108.500 157.000 108.900 ;
        RECT 150.900 107.700 151.300 107.800 ;
        RECT 149.400 107.400 151.300 107.700 ;
        RECT 149.400 105.700 149.800 107.400 ;
        RECT 152.900 107.100 153.300 107.200 ;
        RECT 155.800 107.100 156.100 107.800 ;
        RECT 158.200 107.500 158.600 109.900 ;
        RECT 159.000 108.000 159.400 109.900 ;
        RECT 160.600 108.000 161.000 109.900 ;
        RECT 159.000 107.900 161.000 108.000 ;
        RECT 161.400 107.900 161.800 109.900 ;
        RECT 162.200 108.000 162.600 109.900 ;
        RECT 163.800 109.600 165.800 109.900 ;
        RECT 163.800 108.000 164.200 109.600 ;
        RECT 162.200 107.900 164.200 108.000 ;
        RECT 164.600 107.900 165.000 109.300 ;
        RECT 165.400 107.900 165.800 109.600 ;
        RECT 167.800 107.900 168.200 109.900 ;
        RECT 168.500 108.200 168.900 108.600 ;
        RECT 159.100 107.700 160.900 107.900 ;
        RECT 159.400 107.200 159.800 107.400 ;
        RECT 161.400 107.200 161.700 107.900 ;
        RECT 162.300 107.700 164.100 107.900 ;
        RECT 162.600 107.200 163.000 107.400 ;
        RECT 164.700 107.200 165.000 107.900 ;
        RECT 157.400 107.100 158.200 107.200 ;
        RECT 152.700 106.800 158.200 107.100 ;
        RECT 159.000 106.900 159.800 107.200 ;
        RECT 159.000 106.800 159.400 106.900 ;
        RECT 160.500 106.800 161.800 107.200 ;
        RECT 162.200 106.900 163.000 107.200 ;
        RECT 163.800 106.900 165.000 107.200 ;
        RECT 162.200 106.800 162.600 106.900 ;
        RECT 163.800 106.800 164.200 106.900 ;
        RECT 151.800 106.400 152.200 106.500 ;
        RECT 150.300 106.100 152.200 106.400 ;
        RECT 150.300 106.000 150.700 106.100 ;
        RECT 151.100 105.700 151.500 105.800 ;
        RECT 149.400 105.400 151.500 105.700 ;
        RECT 149.400 101.100 149.800 105.400 ;
        RECT 152.700 105.200 153.000 106.800 ;
        RECT 156.300 106.700 156.700 106.800 ;
        RECT 155.800 106.200 156.200 106.300 ;
        RECT 157.100 106.200 157.500 106.300 ;
        RECT 155.000 105.900 157.500 106.200 ;
        RECT 155.000 105.800 155.400 105.900 ;
        RECT 159.800 105.800 160.200 106.600 ;
        RECT 155.800 105.500 158.600 105.600 ;
        RECT 155.700 105.400 158.600 105.500 ;
        RECT 151.800 104.900 153.000 105.200 ;
        RECT 153.700 105.300 158.600 105.400 ;
        RECT 153.700 105.100 156.100 105.300 ;
        RECT 151.800 104.400 152.100 104.900 ;
        RECT 151.400 104.000 152.100 104.400 ;
        RECT 152.900 104.500 153.300 104.600 ;
        RECT 153.700 104.500 154.000 105.100 ;
        RECT 152.900 104.200 154.000 104.500 ;
        RECT 154.300 104.500 157.000 104.800 ;
        RECT 154.300 104.400 154.700 104.500 ;
        RECT 156.600 104.400 157.000 104.500 ;
        RECT 153.500 103.700 153.900 103.800 ;
        RECT 154.900 103.700 155.300 103.800 ;
        RECT 151.800 103.100 152.200 103.500 ;
        RECT 153.500 103.400 155.300 103.700 ;
        RECT 153.900 103.100 154.200 103.400 ;
        RECT 156.600 103.100 157.000 103.500 ;
        RECT 151.500 101.100 152.100 103.100 ;
        RECT 153.800 101.100 154.200 103.100 ;
        RECT 156.000 102.800 157.000 103.100 ;
        RECT 156.000 101.100 156.400 102.800 ;
        RECT 158.200 101.100 158.600 105.300 ;
        RECT 160.500 105.100 160.800 106.800 ;
        RECT 163.000 105.800 163.400 106.600 ;
        RECT 161.400 105.100 161.800 105.200 ;
        RECT 163.800 105.100 164.100 106.800 ;
        RECT 164.600 105.800 165.000 106.600 ;
        RECT 165.400 106.400 165.800 107.200 ;
        RECT 167.000 106.400 167.400 107.200 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 167.800 106.100 168.100 107.900 ;
        RECT 168.600 107.800 169.000 108.200 ;
        RECT 168.600 106.100 169.000 106.200 ;
        RECT 166.200 105.800 167.000 106.100 ;
        RECT 167.800 105.800 169.000 106.100 ;
        RECT 169.400 106.100 169.800 109.900 ;
        RECT 170.200 108.100 170.600 108.600 ;
        RECT 171.000 108.100 171.400 109.900 ;
        RECT 173.100 109.200 173.700 109.900 ;
        RECT 173.100 108.900 173.800 109.200 ;
        RECT 175.400 108.900 175.800 109.900 ;
        RECT 177.600 109.200 178.000 109.900 ;
        RECT 177.600 108.900 178.600 109.200 ;
        RECT 173.400 108.500 173.800 108.900 ;
        RECT 175.500 108.600 175.800 108.900 ;
        RECT 175.500 108.300 176.900 108.600 ;
        RECT 176.500 108.200 176.900 108.300 ;
        RECT 177.400 108.200 177.800 108.600 ;
        RECT 178.200 108.500 178.600 108.900 ;
        RECT 170.200 107.800 171.400 108.100 ;
        RECT 171.000 107.700 171.400 107.800 ;
        RECT 172.500 107.700 172.900 107.800 ;
        RECT 171.000 107.400 172.900 107.700 ;
        RECT 170.200 106.100 170.600 106.200 ;
        RECT 169.400 105.800 170.600 106.100 ;
        RECT 166.600 105.600 167.000 105.800 ;
        RECT 168.600 105.100 168.900 105.800 ;
        RECT 160.300 104.800 160.800 105.100 ;
        RECT 161.100 104.800 161.800 105.100 ;
        RECT 160.300 101.100 160.700 104.800 ;
        RECT 161.100 104.200 161.400 104.800 ;
        RECT 161.000 103.800 161.400 104.200 ;
        RECT 163.500 101.100 164.500 105.100 ;
        RECT 166.200 104.800 168.200 105.100 ;
        RECT 166.200 101.100 166.600 104.800 ;
        RECT 167.800 101.100 168.200 104.800 ;
        RECT 168.600 101.100 169.000 105.100 ;
        RECT 169.400 101.100 169.800 105.800 ;
        RECT 171.000 105.700 171.400 107.400 ;
        RECT 174.500 107.100 174.900 107.200 ;
        RECT 176.600 107.100 177.000 107.200 ;
        RECT 177.400 107.100 177.700 108.200 ;
        RECT 179.800 107.500 180.200 109.900 ;
        RECT 179.000 107.100 179.800 107.200 ;
        RECT 174.300 106.800 179.800 107.100 ;
        RECT 173.400 106.400 173.800 106.500 ;
        RECT 171.900 106.100 173.800 106.400 ;
        RECT 171.900 106.000 172.300 106.100 ;
        RECT 172.700 105.700 173.100 105.800 ;
        RECT 171.000 105.400 173.100 105.700 ;
        RECT 171.000 101.100 171.400 105.400 ;
        RECT 174.300 105.200 174.600 106.800 ;
        RECT 177.900 106.700 178.300 106.800 ;
        RECT 178.700 106.200 179.100 106.300 ;
        RECT 176.600 105.900 179.100 106.200 ;
        RECT 176.600 105.800 177.000 105.900 ;
        RECT 177.400 105.500 180.200 105.600 ;
        RECT 177.300 105.400 180.200 105.500 ;
        RECT 173.400 104.900 174.600 105.200 ;
        RECT 175.300 105.300 180.200 105.400 ;
        RECT 175.300 105.100 177.700 105.300 ;
        RECT 173.400 104.400 173.700 104.900 ;
        RECT 173.000 104.200 173.700 104.400 ;
        RECT 174.500 104.500 174.900 104.600 ;
        RECT 175.300 104.500 175.600 105.100 ;
        RECT 174.500 104.200 175.600 104.500 ;
        RECT 175.900 104.500 178.600 104.800 ;
        RECT 175.900 104.400 176.300 104.500 ;
        RECT 178.200 104.400 178.600 104.500 ;
        RECT 172.600 104.000 173.700 104.200 ;
        RECT 172.600 103.800 173.300 104.000 ;
        RECT 175.100 103.700 175.500 103.800 ;
        RECT 176.500 103.700 176.900 103.800 ;
        RECT 173.400 103.100 173.800 103.500 ;
        RECT 175.100 103.400 176.900 103.700 ;
        RECT 175.500 103.100 175.800 103.400 ;
        RECT 178.200 103.100 178.600 103.500 ;
        RECT 173.100 101.100 173.700 103.100 ;
        RECT 175.400 101.100 175.800 103.100 ;
        RECT 177.600 102.800 178.600 103.100 ;
        RECT 177.600 101.100 178.000 102.800 ;
        RECT 179.800 101.100 180.200 105.300 ;
        RECT 0.600 95.700 1.000 99.900 ;
        RECT 2.800 98.200 3.200 99.900 ;
        RECT 2.200 97.900 3.200 98.200 ;
        RECT 5.000 97.900 5.400 99.900 ;
        RECT 7.100 97.900 7.700 99.900 ;
        RECT 2.200 97.500 2.600 97.900 ;
        RECT 5.000 97.600 5.300 97.900 ;
        RECT 3.900 97.300 5.700 97.600 ;
        RECT 7.000 97.500 7.400 97.900 ;
        RECT 3.900 97.200 4.300 97.300 ;
        RECT 5.300 97.200 5.700 97.300 ;
        RECT 2.200 96.500 2.600 96.600 ;
        RECT 4.500 96.500 4.900 96.600 ;
        RECT 2.200 96.200 4.900 96.500 ;
        RECT 5.200 96.500 6.300 96.800 ;
        RECT 5.200 95.900 5.500 96.500 ;
        RECT 5.900 96.400 6.300 96.500 ;
        RECT 7.100 96.600 7.800 97.000 ;
        RECT 7.100 96.100 7.400 96.600 ;
        RECT 3.100 95.700 5.500 95.900 ;
        RECT 0.600 95.600 5.500 95.700 ;
        RECT 6.200 95.800 7.400 96.100 ;
        RECT 0.600 95.500 3.500 95.600 ;
        RECT 0.600 95.400 3.400 95.500 ;
        RECT 3.800 95.100 4.200 95.200 ;
        RECT 1.700 94.800 4.200 95.100 ;
        RECT 1.700 94.700 2.100 94.800 ;
        RECT 2.500 94.200 2.900 94.300 ;
        RECT 6.200 94.200 6.500 95.800 ;
        RECT 9.400 95.600 9.800 99.900 ;
        RECT 7.700 95.300 9.800 95.600 ;
        RECT 7.700 95.200 8.100 95.300 ;
        RECT 8.500 94.900 8.900 95.000 ;
        RECT 7.000 94.600 8.900 94.900 ;
        RECT 7.000 94.500 7.400 94.600 ;
        RECT 1.000 93.900 6.500 94.200 ;
        RECT 1.000 93.800 1.800 93.900 ;
        RECT 0.600 91.100 1.000 93.500 ;
        RECT 3.100 93.200 3.400 93.900 ;
        RECT 5.900 93.800 6.300 93.900 ;
        RECT 9.400 93.600 9.800 95.300 ;
        RECT 7.900 93.300 9.800 93.600 ;
        RECT 7.900 93.200 8.300 93.300 ;
        RECT 2.200 92.100 2.600 92.500 ;
        RECT 3.000 92.400 3.400 93.200 ;
        RECT 9.400 93.100 9.800 93.300 ;
        RECT 11.000 95.100 11.400 99.900 ;
        RECT 13.700 96.400 14.100 99.900 ;
        RECT 15.800 97.500 16.200 99.500 ;
        RECT 13.300 96.100 14.100 96.400 ;
        RECT 12.600 95.100 13.000 95.600 ;
        RECT 11.000 94.800 13.000 95.100 ;
        RECT 10.200 93.100 10.600 93.200 ;
        RECT 9.400 92.800 10.600 93.100 ;
        RECT 3.900 92.700 4.300 92.800 ;
        RECT 3.900 92.400 5.300 92.700 ;
        RECT 5.000 92.100 5.300 92.400 ;
        RECT 7.000 92.100 7.400 92.500 ;
        RECT 2.200 91.800 3.200 92.100 ;
        RECT 2.800 91.100 3.200 91.800 ;
        RECT 5.000 91.100 5.400 92.100 ;
        RECT 7.000 91.800 7.700 92.100 ;
        RECT 7.100 91.100 7.700 91.800 ;
        RECT 9.400 91.100 9.800 92.800 ;
        RECT 10.200 92.400 10.600 92.800 ;
        RECT 11.000 91.100 11.400 94.800 ;
        RECT 13.300 94.200 13.600 96.100 ;
        RECT 15.900 95.800 16.200 97.500 ;
        RECT 16.600 96.200 17.000 99.900 ;
        RECT 18.200 99.600 20.200 99.900 ;
        RECT 18.200 96.200 18.600 99.600 ;
        RECT 16.600 95.900 18.600 96.200 ;
        RECT 19.000 95.900 19.400 99.300 ;
        RECT 19.800 95.900 20.200 99.600 ;
        RECT 20.900 96.300 21.300 99.900 ;
        RECT 20.900 95.900 21.800 96.300 ;
        RECT 23.000 95.900 23.400 99.900 ;
        RECT 23.800 96.200 24.200 99.900 ;
        RECT 25.400 96.200 25.800 99.900 ;
        RECT 23.800 95.900 25.800 96.200 ;
        RECT 14.300 95.500 16.200 95.800 ;
        RECT 19.000 95.600 19.300 95.900 ;
        RECT 14.300 94.500 14.600 95.500 ;
        RECT 17.000 95.200 17.400 95.400 ;
        RECT 18.300 95.300 19.300 95.600 ;
        RECT 18.300 95.200 18.600 95.300 ;
        RECT 11.800 94.100 12.200 94.200 ;
        RECT 12.600 94.100 13.600 94.200 ;
        RECT 13.900 94.100 14.600 94.500 ;
        RECT 15.000 94.400 15.400 95.200 ;
        RECT 15.800 94.400 16.200 95.200 ;
        RECT 16.600 94.900 17.400 95.200 ;
        RECT 16.600 94.800 17.000 94.900 ;
        RECT 18.200 94.800 18.600 95.200 ;
        RECT 19.800 94.800 20.200 95.600 ;
        RECT 20.600 94.800 21.000 95.600 ;
        RECT 11.800 93.800 13.600 94.100 ;
        RECT 13.300 93.500 13.600 93.800 ;
        RECT 14.100 93.900 14.600 94.100 ;
        RECT 14.100 93.600 16.200 93.900 ;
        RECT 17.400 93.800 17.800 94.600 ;
        RECT 13.300 93.300 13.700 93.500 ;
        RECT 13.300 93.000 14.100 93.300 ;
        RECT 13.700 91.500 14.100 93.000 ;
        RECT 15.900 92.500 16.200 93.600 ;
        RECT 18.300 93.100 18.600 94.800 ;
        RECT 18.900 94.400 19.300 94.800 ;
        RECT 19.000 94.200 19.300 94.400 ;
        RECT 21.400 94.200 21.700 95.900 ;
        RECT 23.100 95.200 23.400 95.900 ;
        RECT 26.200 95.600 26.600 99.900 ;
        RECT 28.300 97.900 28.900 99.900 ;
        RECT 30.600 97.900 31.000 99.900 ;
        RECT 32.800 98.200 33.200 99.900 ;
        RECT 32.800 97.900 33.800 98.200 ;
        RECT 28.600 97.500 29.000 97.900 ;
        RECT 30.700 97.600 31.000 97.900 ;
        RECT 30.300 97.300 32.100 97.600 ;
        RECT 33.400 97.500 33.800 97.900 ;
        RECT 30.300 97.200 30.700 97.300 ;
        RECT 31.700 97.200 32.100 97.300 ;
        RECT 28.200 96.600 28.900 97.000 ;
        RECT 28.600 96.100 28.900 96.600 ;
        RECT 29.700 96.500 30.800 96.800 ;
        RECT 29.700 96.400 30.100 96.500 ;
        RECT 28.600 95.800 29.800 96.100 ;
        RECT 25.000 95.200 25.400 95.400 ;
        RECT 26.200 95.300 28.300 95.600 ;
        RECT 23.000 94.900 24.200 95.200 ;
        RECT 25.000 94.900 25.800 95.200 ;
        RECT 23.000 94.800 23.400 94.900 ;
        RECT 23.800 94.800 24.200 94.900 ;
        RECT 25.400 94.800 25.800 94.900 ;
        RECT 19.000 94.100 19.400 94.200 ;
        RECT 20.600 94.100 21.000 94.200 ;
        RECT 19.000 93.800 21.000 94.100 ;
        RECT 21.400 94.100 21.800 94.200 ;
        RECT 21.400 93.800 23.300 94.100 ;
        RECT 15.800 91.500 16.200 92.500 ;
        RECT 18.100 92.200 18.900 93.100 ;
        RECT 18.100 91.800 19.400 92.200 ;
        RECT 21.400 92.100 21.700 93.800 ;
        RECT 23.000 93.200 23.300 93.800 ;
        RECT 22.200 92.400 22.600 93.200 ;
        RECT 23.000 92.800 23.400 93.200 ;
        RECT 23.900 93.100 24.200 94.800 ;
        RECT 24.600 93.800 25.000 94.600 ;
        RECT 23.100 92.400 23.500 92.800 ;
        RECT 18.100 91.100 18.900 91.800 ;
        RECT 21.400 91.100 21.800 92.100 ;
        RECT 23.800 91.100 24.200 93.100 ;
        RECT 26.200 93.600 26.600 95.300 ;
        RECT 27.900 95.200 28.300 95.300 ;
        RECT 27.100 94.900 27.500 95.000 ;
        RECT 27.100 94.600 29.000 94.900 ;
        RECT 28.600 94.500 29.000 94.600 ;
        RECT 29.500 94.200 29.800 95.800 ;
        RECT 30.500 95.900 30.800 96.500 ;
        RECT 31.100 96.500 31.500 96.600 ;
        RECT 33.400 96.500 33.800 96.600 ;
        RECT 31.100 96.200 33.800 96.500 ;
        RECT 30.500 95.700 32.900 95.900 ;
        RECT 35.000 95.700 35.400 99.900 ;
        RECT 36.600 97.900 37.000 99.900 ;
        RECT 36.700 97.800 37.000 97.900 ;
        RECT 38.200 97.900 38.600 99.900 ;
        RECT 41.400 97.900 41.800 99.900 ;
        RECT 38.200 97.800 38.500 97.900 ;
        RECT 36.700 97.500 38.500 97.800 ;
        RECT 37.400 96.400 37.800 97.200 ;
        RECT 38.200 96.200 38.500 97.500 ;
        RECT 30.500 95.600 35.400 95.700 ;
        RECT 32.500 95.500 35.400 95.600 ;
        RECT 32.600 95.400 35.400 95.500 ;
        RECT 35.800 95.400 36.200 96.200 ;
        RECT 38.200 95.800 38.600 96.200 ;
        RECT 41.500 95.800 41.800 97.900 ;
        RECT 43.000 95.900 43.400 99.900 ;
        RECT 43.800 97.900 44.200 99.900 ;
        RECT 43.900 97.800 44.200 97.900 ;
        RECT 45.400 97.900 45.800 99.900 ;
        RECT 47.800 97.900 48.200 99.900 ;
        RECT 45.400 97.800 45.700 97.900 ;
        RECT 43.900 97.500 45.700 97.800 ;
        RECT 47.900 97.800 48.200 97.900 ;
        RECT 49.400 97.900 49.800 99.900 ;
        RECT 49.400 97.800 49.700 97.900 ;
        RECT 47.900 97.500 49.700 97.800 ;
        RECT 43.900 96.200 44.200 97.500 ;
        RECT 44.600 96.400 45.000 97.200 ;
        RECT 48.600 96.400 49.000 97.200 ;
        RECT 49.400 96.200 49.700 97.500 ;
        RECT 30.200 95.100 30.600 95.200 ;
        RECT 31.800 95.100 32.200 95.200 ;
        RECT 30.200 94.800 34.300 95.100 ;
        RECT 36.600 94.800 37.400 95.200 ;
        RECT 33.900 94.700 34.300 94.800 ;
        RECT 33.100 94.200 33.500 94.300 ;
        RECT 38.200 94.200 38.500 95.800 ;
        RECT 41.500 95.500 42.700 95.800 ;
        RECT 41.400 94.800 41.800 95.200 ;
        RECT 29.500 93.900 35.000 94.200 ;
        RECT 37.700 94.100 38.500 94.200 ;
        RECT 29.700 93.800 30.100 93.900 ;
        RECT 31.000 93.800 31.400 93.900 ;
        RECT 26.200 93.300 28.100 93.600 ;
        RECT 26.200 91.100 26.600 93.300 ;
        RECT 27.700 93.200 28.100 93.300 ;
        RECT 32.600 92.800 32.900 93.900 ;
        RECT 34.200 93.800 35.000 93.900 ;
        RECT 37.600 93.900 38.500 94.100 ;
        RECT 31.700 92.700 32.100 92.800 ;
        RECT 28.600 92.100 29.000 92.500 ;
        RECT 30.700 92.400 32.100 92.700 ;
        RECT 32.600 92.400 33.000 92.800 ;
        RECT 30.700 92.100 31.000 92.400 ;
        RECT 33.400 92.100 33.800 92.500 ;
        RECT 28.300 91.800 29.000 92.100 ;
        RECT 28.300 91.100 28.900 91.800 ;
        RECT 30.600 91.100 31.000 92.100 ;
        RECT 32.800 91.800 33.800 92.100 ;
        RECT 32.800 91.100 33.200 91.800 ;
        RECT 35.000 91.100 35.400 93.500 ;
        RECT 36.600 92.100 37.000 92.200 ;
        RECT 37.600 92.100 38.000 93.900 ;
        RECT 40.600 93.800 41.000 94.600 ;
        RECT 41.500 94.400 41.800 94.800 ;
        RECT 41.500 94.100 42.000 94.400 ;
        RECT 41.600 94.000 42.000 94.100 ;
        RECT 42.400 93.800 42.700 95.500 ;
        RECT 43.100 95.200 43.400 95.900 ;
        RECT 43.800 95.800 44.200 96.200 ;
        RECT 43.000 94.800 43.400 95.200 ;
        RECT 42.400 93.700 42.800 93.800 ;
        RECT 41.300 93.500 42.800 93.700 ;
        RECT 40.700 93.400 42.800 93.500 ;
        RECT 40.700 93.200 41.600 93.400 ;
        RECT 40.700 93.100 41.000 93.200 ;
        RECT 43.100 93.100 43.400 94.800 ;
        RECT 43.900 94.200 44.200 95.800 ;
        RECT 46.200 95.400 46.600 96.200 ;
        RECT 47.000 95.400 47.400 96.200 ;
        RECT 49.400 95.800 49.800 96.200 ;
        RECT 50.200 95.800 50.600 96.600 ;
        RECT 45.000 94.800 45.800 95.200 ;
        RECT 47.800 94.800 48.600 95.200 ;
        RECT 49.400 94.200 49.700 95.800 ;
        RECT 43.900 94.100 44.700 94.200 ;
        RECT 48.900 94.100 49.700 94.200 ;
        RECT 43.900 93.900 44.800 94.100 ;
        RECT 36.600 91.800 38.000 92.100 ;
        RECT 37.600 91.100 38.000 91.800 ;
        RECT 40.600 91.100 41.000 93.100 ;
        RECT 42.700 92.600 43.400 93.100 ;
        RECT 42.700 92.200 43.100 92.600 ;
        RECT 42.700 91.800 43.400 92.200 ;
        RECT 42.700 91.100 43.100 91.800 ;
        RECT 44.400 91.100 44.800 93.900 ;
        RECT 48.800 93.900 49.700 94.100 ;
        RECT 48.800 91.100 49.200 93.900 ;
        RECT 51.000 93.100 51.400 99.900 ;
        RECT 52.700 99.600 54.500 99.900 ;
        RECT 52.700 99.500 53.000 99.600 ;
        RECT 52.600 96.500 53.000 99.500 ;
        RECT 54.200 99.500 54.500 99.600 ;
        RECT 55.000 99.600 57.000 99.900 ;
        RECT 53.400 96.500 53.800 99.300 ;
        RECT 54.200 96.700 54.600 99.500 ;
        RECT 55.000 97.000 55.400 99.600 ;
        RECT 55.800 96.900 56.200 99.300 ;
        RECT 56.600 96.900 57.000 99.600 ;
        RECT 55.800 96.700 56.100 96.900 ;
        RECT 54.200 96.500 56.100 96.700 ;
        RECT 53.500 96.200 53.800 96.500 ;
        RECT 54.300 96.400 56.100 96.500 ;
        RECT 56.700 96.600 57.000 96.900 ;
        RECT 58.200 96.900 58.600 99.900 ;
        RECT 58.200 96.600 58.500 96.900 ;
        RECT 56.700 96.300 58.500 96.600 ;
        RECT 53.400 96.100 53.800 96.200 ;
        RECT 53.400 95.800 55.100 96.100 ;
        RECT 51.800 93.400 52.200 94.200 ;
        RECT 50.500 92.800 51.400 93.100 ;
        RECT 50.500 91.100 50.900 92.800 ;
        RECT 54.800 92.500 55.100 95.800 ;
        RECT 59.000 95.700 59.400 99.900 ;
        RECT 61.200 98.200 61.600 99.900 ;
        RECT 60.600 97.900 61.600 98.200 ;
        RECT 63.400 97.900 63.800 99.900 ;
        RECT 65.500 97.900 66.100 99.900 ;
        RECT 60.600 97.500 61.000 97.900 ;
        RECT 63.400 97.600 63.700 97.900 ;
        RECT 62.300 97.300 64.100 97.600 ;
        RECT 65.400 97.500 65.800 97.900 ;
        RECT 62.300 97.200 62.700 97.300 ;
        RECT 63.700 97.200 64.100 97.300 ;
        RECT 60.600 96.500 61.000 96.600 ;
        RECT 62.900 96.500 63.300 96.600 ;
        RECT 60.600 96.200 63.300 96.500 ;
        RECT 63.600 96.500 64.700 96.800 ;
        RECT 63.600 95.900 63.900 96.500 ;
        RECT 64.300 96.400 64.700 96.500 ;
        RECT 65.500 96.600 66.200 97.000 ;
        RECT 65.500 96.100 65.800 96.600 ;
        RECT 61.500 95.700 63.900 95.900 ;
        RECT 59.000 95.600 63.900 95.700 ;
        RECT 64.600 95.800 65.800 96.100 ;
        RECT 59.000 95.500 61.900 95.600 ;
        RECT 59.000 95.400 61.800 95.500 ;
        RECT 64.600 95.200 64.900 95.800 ;
        RECT 67.800 95.600 68.200 99.900 ;
        RECT 66.100 95.300 68.200 95.600 ;
        RECT 66.100 95.200 66.500 95.300 ;
        RECT 55.400 95.100 56.200 95.200 ;
        RECT 57.400 95.100 57.800 95.200 ;
        RECT 62.200 95.100 62.600 95.200 ;
        RECT 55.400 94.800 57.800 95.100 ;
        RECT 60.100 94.800 62.600 95.100 ;
        RECT 64.600 94.800 65.000 95.200 ;
        RECT 66.900 94.900 67.300 95.000 ;
        RECT 60.100 94.700 60.500 94.800 ;
        RECT 60.900 94.200 61.300 94.300 ;
        RECT 64.600 94.200 64.900 94.800 ;
        RECT 65.400 94.600 67.300 94.900 ;
        RECT 65.400 94.500 65.800 94.600 ;
        RECT 56.200 93.800 57.000 94.200 ;
        RECT 59.400 93.900 64.900 94.200 ;
        RECT 59.400 93.800 60.200 93.900 ;
        RECT 56.900 92.800 57.800 93.200 ;
        RECT 54.800 92.200 56.800 92.500 ;
        RECT 54.800 92.100 55.400 92.200 ;
        RECT 55.000 91.100 55.400 92.100 ;
        RECT 56.500 91.800 57.000 92.200 ;
        RECT 56.600 91.100 57.000 91.800 ;
        RECT 59.000 91.100 59.400 93.500 ;
        RECT 61.500 92.800 61.800 93.900 ;
        RECT 64.300 93.800 64.700 93.900 ;
        RECT 67.800 93.600 68.200 95.300 ;
        RECT 66.300 93.300 68.200 93.600 ;
        RECT 66.300 93.200 66.700 93.300 ;
        RECT 67.800 93.100 68.200 93.300 ;
        RECT 69.400 95.100 69.800 99.900 ;
        RECT 72.100 96.400 72.500 99.900 ;
        RECT 74.200 97.500 74.600 99.500 ;
        RECT 71.700 96.100 72.500 96.400 ;
        RECT 71.000 95.100 71.400 95.600 ;
        RECT 69.400 94.800 71.400 95.100 ;
        RECT 68.600 93.100 69.000 93.200 ;
        RECT 67.800 92.800 69.000 93.100 ;
        RECT 60.600 92.100 61.000 92.500 ;
        RECT 61.400 92.400 61.800 92.800 ;
        RECT 62.300 92.700 62.700 92.800 ;
        RECT 62.300 92.400 63.700 92.700 ;
        RECT 63.400 92.100 63.700 92.400 ;
        RECT 65.400 92.100 65.800 92.500 ;
        RECT 60.600 91.800 61.600 92.100 ;
        RECT 61.200 91.100 61.600 91.800 ;
        RECT 63.400 91.100 63.800 92.100 ;
        RECT 65.400 91.800 66.100 92.100 ;
        RECT 65.500 91.100 66.100 91.800 ;
        RECT 67.800 91.100 68.200 92.800 ;
        RECT 68.600 92.400 69.000 92.800 ;
        RECT 69.400 91.100 69.800 94.800 ;
        RECT 71.700 94.200 72.000 96.100 ;
        RECT 74.300 95.800 74.600 97.500 ;
        RECT 72.700 95.500 74.600 95.800 ;
        RECT 75.000 95.600 75.400 99.900 ;
        RECT 77.100 97.900 77.700 99.900 ;
        RECT 79.400 97.900 79.800 99.900 ;
        RECT 81.600 98.200 82.000 99.900 ;
        RECT 81.600 97.900 82.600 98.200 ;
        RECT 77.400 97.500 77.800 97.900 ;
        RECT 79.500 97.600 79.800 97.900 ;
        RECT 79.100 97.300 80.900 97.600 ;
        RECT 82.200 97.500 82.600 97.900 ;
        RECT 79.100 97.200 79.500 97.300 ;
        RECT 80.500 97.200 80.900 97.300 ;
        RECT 76.600 97.000 77.300 97.200 ;
        RECT 76.600 96.800 77.700 97.000 ;
        RECT 77.000 96.600 77.700 96.800 ;
        RECT 77.400 96.100 77.700 96.600 ;
        RECT 78.500 96.500 79.600 96.800 ;
        RECT 78.500 96.400 78.900 96.500 ;
        RECT 77.400 95.800 78.600 96.100 ;
        RECT 72.700 94.500 73.000 95.500 ;
        RECT 75.000 95.300 77.100 95.600 ;
        RECT 70.200 94.100 70.600 94.200 ;
        RECT 71.000 94.100 72.000 94.200 ;
        RECT 72.300 94.100 73.000 94.500 ;
        RECT 73.400 94.400 73.800 95.200 ;
        RECT 74.200 94.400 74.600 95.200 ;
        RECT 70.200 93.800 72.000 94.100 ;
        RECT 71.700 93.500 72.000 93.800 ;
        RECT 72.500 93.900 73.000 94.100 ;
        RECT 72.500 93.600 74.600 93.900 ;
        RECT 71.700 93.300 72.100 93.500 ;
        RECT 71.700 93.000 72.500 93.300 ;
        RECT 72.100 91.500 72.500 93.000 ;
        RECT 74.300 92.500 74.600 93.600 ;
        RECT 74.200 91.500 74.600 92.500 ;
        RECT 75.000 93.600 75.400 95.300 ;
        RECT 76.700 95.200 77.100 95.300 ;
        RECT 75.900 94.900 76.300 95.000 ;
        RECT 75.900 94.600 77.800 94.900 ;
        RECT 77.400 94.500 77.800 94.600 ;
        RECT 78.300 94.200 78.600 95.800 ;
        RECT 79.300 95.900 79.600 96.500 ;
        RECT 79.900 96.500 80.300 96.600 ;
        RECT 82.200 96.500 82.600 96.600 ;
        RECT 79.900 96.200 82.600 96.500 ;
        RECT 79.300 95.700 81.700 95.900 ;
        RECT 83.800 95.700 84.200 99.900 ;
        RECT 79.300 95.600 84.200 95.700 ;
        RECT 81.300 95.500 84.200 95.600 ;
        RECT 81.400 95.400 84.200 95.500 ;
        RECT 86.200 95.600 86.600 99.900 ;
        RECT 88.300 97.900 88.900 99.900 ;
        RECT 90.600 97.900 91.000 99.900 ;
        RECT 92.800 98.200 93.200 99.900 ;
        RECT 92.800 97.900 93.800 98.200 ;
        RECT 88.600 97.500 89.000 97.900 ;
        RECT 90.700 97.600 91.000 97.900 ;
        RECT 90.300 97.300 92.100 97.600 ;
        RECT 93.400 97.500 93.800 97.900 ;
        RECT 90.300 97.200 90.700 97.300 ;
        RECT 91.700 97.200 92.100 97.300 ;
        RECT 88.200 96.600 88.900 97.000 ;
        RECT 88.600 96.100 88.900 96.600 ;
        RECT 89.700 96.500 90.800 96.800 ;
        RECT 89.700 96.400 90.100 96.500 ;
        RECT 88.600 95.800 89.800 96.100 ;
        RECT 86.200 95.300 88.300 95.600 ;
        RECT 80.600 95.100 81.000 95.200 ;
        RECT 80.600 94.800 83.100 95.100 ;
        RECT 82.700 94.700 83.100 94.800 ;
        RECT 81.900 94.200 82.300 94.300 ;
        RECT 78.300 93.900 83.800 94.200 ;
        RECT 78.500 93.800 78.900 93.900 ;
        RECT 75.000 93.300 76.900 93.600 ;
        RECT 75.000 91.100 75.400 93.300 ;
        RECT 76.500 93.200 76.900 93.300 ;
        RECT 81.400 92.800 81.700 93.900 ;
        RECT 83.000 93.800 83.800 93.900 ;
        RECT 86.200 93.600 86.600 95.300 ;
        RECT 87.900 95.200 88.300 95.300 ;
        RECT 87.100 94.900 87.500 95.000 ;
        RECT 87.100 94.600 89.000 94.900 ;
        RECT 88.600 94.500 89.000 94.600 ;
        RECT 89.500 94.200 89.800 95.800 ;
        RECT 90.500 95.900 90.800 96.500 ;
        RECT 91.100 96.500 91.500 96.600 ;
        RECT 93.400 96.500 93.800 96.600 ;
        RECT 91.100 96.200 93.800 96.500 ;
        RECT 90.500 95.700 92.900 95.900 ;
        RECT 95.000 95.700 95.400 99.900 ;
        RECT 90.500 95.600 95.400 95.700 ;
        RECT 92.500 95.500 95.400 95.600 ;
        RECT 92.600 95.400 95.400 95.500 ;
        RECT 91.000 95.100 91.400 95.200 ;
        RECT 91.800 95.100 92.200 95.200 ;
        RECT 91.000 94.800 94.300 95.100 ;
        RECT 93.900 94.700 94.300 94.800 ;
        RECT 93.100 94.200 93.500 94.300 ;
        RECT 89.500 93.900 95.000 94.200 ;
        RECT 89.700 93.800 90.100 93.900 ;
        RECT 92.600 93.800 93.000 93.900 ;
        RECT 94.200 93.800 95.000 93.900 ;
        RECT 80.500 92.700 80.900 92.800 ;
        RECT 77.400 92.100 77.800 92.500 ;
        RECT 79.500 92.400 80.900 92.700 ;
        RECT 81.400 92.400 81.800 92.800 ;
        RECT 79.500 92.100 79.800 92.400 ;
        RECT 82.200 92.100 82.600 92.500 ;
        RECT 77.100 91.800 77.800 92.100 ;
        RECT 77.100 91.100 77.700 91.800 ;
        RECT 79.400 91.100 79.800 92.100 ;
        RECT 81.600 91.800 82.600 92.100 ;
        RECT 81.600 91.100 82.000 91.800 ;
        RECT 83.800 91.100 84.200 93.500 ;
        RECT 86.200 93.300 88.100 93.600 ;
        RECT 85.400 92.100 85.800 92.200 ;
        RECT 86.200 92.100 86.600 93.300 ;
        RECT 87.700 93.200 88.100 93.300 ;
        RECT 92.600 92.800 92.900 93.800 ;
        RECT 91.700 92.700 92.100 92.800 ;
        RECT 88.600 92.100 89.000 92.500 ;
        RECT 90.700 92.400 92.100 92.700 ;
        RECT 92.600 92.400 93.000 92.800 ;
        RECT 90.700 92.100 91.000 92.400 ;
        RECT 93.400 92.100 93.800 92.500 ;
        RECT 85.400 91.800 86.600 92.100 ;
        RECT 86.200 91.100 86.600 91.800 ;
        RECT 88.300 91.800 89.000 92.100 ;
        RECT 88.300 91.100 88.900 91.800 ;
        RECT 90.600 91.100 91.000 92.100 ;
        RECT 92.800 91.800 93.800 92.100 ;
        RECT 92.800 91.100 93.200 91.800 ;
        RECT 95.000 91.100 95.400 93.500 ;
        RECT 95.800 93.400 96.200 94.200 ;
        RECT 96.600 93.100 97.000 99.900 ;
        RECT 97.400 95.800 97.800 96.600 ;
        RECT 98.200 93.400 98.600 94.200 ;
        RECT 99.000 93.100 99.400 99.900 ;
        RECT 99.800 95.800 100.200 96.600 ;
        RECT 100.600 95.600 101.000 99.900 ;
        RECT 102.700 97.900 103.300 99.900 ;
        RECT 105.000 97.900 105.400 99.900 ;
        RECT 107.200 98.200 107.600 99.900 ;
        RECT 107.200 97.900 108.200 98.200 ;
        RECT 103.000 97.500 103.400 97.900 ;
        RECT 105.100 97.600 105.400 97.900 ;
        RECT 104.700 97.300 106.500 97.600 ;
        RECT 107.800 97.500 108.200 97.900 ;
        RECT 104.700 97.200 105.100 97.300 ;
        RECT 106.100 97.200 106.500 97.300 ;
        RECT 102.600 96.600 103.300 97.000 ;
        RECT 103.000 96.100 103.300 96.600 ;
        RECT 104.100 96.500 105.200 96.800 ;
        RECT 104.100 96.400 104.500 96.500 ;
        RECT 103.000 95.800 104.200 96.100 ;
        RECT 100.600 95.300 102.700 95.600 ;
        RECT 100.600 93.600 101.000 95.300 ;
        RECT 102.300 95.200 102.700 95.300 ;
        RECT 101.500 94.900 101.900 95.000 ;
        RECT 101.500 94.600 103.400 94.900 ;
        RECT 103.000 94.500 103.400 94.600 ;
        RECT 103.900 94.200 104.200 95.800 ;
        RECT 104.900 95.900 105.200 96.500 ;
        RECT 105.500 96.500 105.900 96.600 ;
        RECT 107.800 96.500 108.200 96.600 ;
        RECT 105.500 96.200 108.200 96.500 ;
        RECT 104.900 95.700 107.300 95.900 ;
        RECT 109.400 95.700 109.800 99.900 ;
        RECT 112.100 99.200 112.500 99.900 ;
        RECT 112.100 98.800 113.000 99.200 ;
        RECT 112.100 96.400 112.500 98.800 ;
        RECT 114.200 97.500 114.600 99.500 ;
        RECT 104.900 95.600 109.800 95.700 ;
        RECT 111.700 96.100 112.500 96.400 ;
        RECT 106.900 95.500 109.800 95.600 ;
        RECT 107.000 95.400 109.800 95.500 ;
        RECT 104.600 95.100 105.000 95.200 ;
        RECT 106.200 95.100 106.600 95.200 ;
        RECT 110.200 95.100 110.600 95.200 ;
        RECT 111.000 95.100 111.400 95.600 ;
        RECT 104.600 94.800 108.700 95.100 ;
        RECT 110.200 94.800 111.400 95.100 ;
        RECT 108.300 94.700 108.700 94.800 ;
        RECT 107.500 94.200 107.900 94.300 ;
        RECT 111.700 94.200 112.000 96.100 ;
        RECT 114.300 95.800 114.600 97.500 ;
        RECT 115.300 96.300 115.700 99.900 ;
        RECT 115.300 95.900 116.200 96.300 ;
        RECT 118.200 96.000 118.600 99.900 ;
        RECT 119.800 97.600 120.200 99.900 ;
        RECT 112.700 95.500 114.600 95.800 ;
        RECT 112.700 94.500 113.000 95.500 ;
        RECT 103.900 93.900 109.400 94.200 ;
        RECT 104.100 93.800 104.500 93.900 ;
        RECT 105.400 93.800 105.800 93.900 ;
        RECT 106.200 93.800 106.600 93.900 ;
        RECT 100.600 93.300 102.500 93.600 ;
        RECT 96.600 92.800 97.500 93.100 ;
        RECT 99.000 92.800 99.900 93.100 ;
        RECT 97.100 91.100 97.500 92.800 ;
        RECT 99.500 92.200 99.900 92.800 ;
        RECT 99.500 91.800 100.200 92.200 ;
        RECT 99.500 91.100 99.900 91.800 ;
        RECT 100.600 91.100 101.000 93.300 ;
        RECT 102.100 93.200 102.500 93.300 ;
        RECT 107.000 92.800 107.300 93.900 ;
        RECT 108.600 93.800 109.400 93.900 ;
        RECT 111.000 93.800 112.000 94.200 ;
        RECT 112.300 94.100 113.000 94.500 ;
        RECT 113.400 94.400 113.800 95.200 ;
        RECT 114.200 94.400 114.600 95.200 ;
        RECT 115.000 94.800 115.400 95.600 ;
        RECT 111.700 93.500 112.000 93.800 ;
        RECT 112.500 93.900 113.000 94.100 ;
        RECT 115.800 94.200 116.100 95.900 ;
        RECT 118.100 95.600 118.600 96.000 ;
        RECT 118.900 97.300 120.200 97.600 ;
        RECT 118.900 96.500 119.200 97.300 ;
        RECT 121.400 97.200 121.800 99.900 ;
        RECT 123.000 98.500 123.400 99.900 ;
        RECT 123.800 98.500 124.200 99.900 ;
        RECT 124.600 98.500 125.000 99.900 ;
        RECT 122.100 97.200 124.200 97.600 ;
        RECT 120.500 96.800 121.800 97.200 ;
        RECT 125.400 96.800 125.800 99.900 ;
        RECT 127.000 97.500 127.400 99.900 ;
        RECT 128.600 97.500 129.000 99.900 ;
        RECT 129.400 98.500 129.800 99.900 ;
        RECT 130.200 98.500 130.600 99.900 ;
        RECT 131.800 97.600 132.200 99.900 ;
        RECT 133.400 98.200 133.800 99.900 ;
        RECT 137.400 98.200 137.800 99.900 ;
        RECT 133.400 97.900 133.900 98.200 ;
        RECT 133.600 97.600 133.900 97.900 ;
        RECT 137.300 97.900 137.800 98.200 ;
        RECT 137.300 97.600 137.600 97.900 ;
        RECT 139.000 97.600 139.400 99.900 ;
        RECT 140.600 98.500 141.000 99.900 ;
        RECT 141.400 98.500 141.800 99.900 ;
        RECT 131.200 97.200 133.300 97.600 ;
        RECT 133.600 97.300 134.600 97.600 ;
        RECT 127.000 96.800 128.300 97.200 ;
        RECT 128.600 96.900 131.500 97.200 ;
        RECT 133.000 97.000 133.300 97.200 ;
        RECT 123.000 96.500 123.400 96.600 ;
        RECT 118.900 96.200 123.400 96.500 ;
        RECT 124.600 96.500 125.000 96.600 ;
        RECT 128.600 96.500 128.900 96.900 ;
        RECT 131.800 96.600 132.500 96.900 ;
        RECT 133.000 96.600 133.800 97.000 ;
        RECT 124.600 96.200 128.900 96.500 ;
        RECT 129.400 96.500 132.500 96.600 ;
        RECT 129.400 96.300 132.100 96.500 ;
        RECT 129.400 96.200 129.800 96.300 ;
        RECT 112.500 93.600 114.600 93.900 ;
        RECT 106.100 92.700 106.500 92.800 ;
        RECT 103.000 92.100 103.400 92.500 ;
        RECT 105.100 92.400 106.500 92.700 ;
        RECT 107.000 92.400 107.400 92.800 ;
        RECT 105.100 92.100 105.400 92.400 ;
        RECT 107.800 92.100 108.200 92.500 ;
        RECT 102.700 91.800 103.400 92.100 ;
        RECT 102.700 91.100 103.300 91.800 ;
        RECT 105.000 91.100 105.400 92.100 ;
        RECT 107.200 91.800 108.200 92.100 ;
        RECT 107.200 91.100 107.600 91.800 ;
        RECT 109.400 91.100 109.800 93.500 ;
        RECT 111.700 93.300 112.100 93.500 ;
        RECT 111.700 93.000 112.500 93.300 ;
        RECT 112.100 91.500 112.500 93.000 ;
        RECT 114.300 92.500 114.600 93.600 ;
        RECT 115.800 93.800 116.200 94.200 ;
        RECT 115.000 93.100 115.400 93.200 ;
        RECT 115.800 93.100 116.100 93.800 ;
        RECT 118.100 93.400 118.500 95.600 ;
        RECT 118.900 95.300 119.200 96.200 ;
        RECT 118.800 95.000 119.200 95.300 ;
        RECT 118.800 94.000 119.100 95.000 ;
        RECT 119.400 94.300 121.300 94.700 ;
        RECT 118.800 93.700 119.400 94.000 ;
        RECT 115.000 92.800 116.100 93.100 ;
        RECT 114.200 91.500 114.600 92.500 ;
        RECT 115.800 92.100 116.100 92.800 ;
        RECT 116.600 93.100 117.000 93.200 ;
        RECT 118.100 93.100 118.600 93.400 ;
        RECT 116.600 92.800 118.600 93.100 ;
        RECT 116.600 92.400 117.000 92.800 ;
        RECT 115.800 91.100 116.200 92.100 ;
        RECT 118.200 91.100 118.600 92.800 ;
        RECT 119.000 91.100 119.400 93.700 ;
        RECT 120.900 93.700 121.300 94.300 ;
        RECT 120.900 93.400 121.800 93.700 ;
        RECT 121.400 93.100 121.800 93.400 ;
        RECT 123.800 93.200 124.200 94.600 ;
        RECT 125.400 94.300 127.000 94.700 ;
        RECT 128.900 94.300 129.900 94.700 ;
        RECT 134.200 94.500 134.600 97.300 ;
        RECT 125.200 93.900 125.600 94.000 ;
        RECT 125.200 93.600 127.400 93.900 ;
        RECT 127.000 93.500 127.400 93.600 ;
        RECT 127.800 93.400 128.200 94.200 ;
        RECT 121.400 92.700 122.600 93.100 ;
        RECT 123.800 92.800 124.300 93.200 ;
        RECT 125.800 92.800 126.600 93.200 ;
        RECT 127.000 93.100 127.400 93.200 ;
        RECT 128.900 93.100 129.300 94.300 ;
        RECT 130.200 94.100 134.600 94.500 ;
        RECT 131.900 93.400 133.400 93.800 ;
        RECT 131.900 93.100 132.300 93.400 ;
        RECT 127.000 92.800 129.300 93.100 ;
        RECT 122.200 91.100 122.600 92.700 ;
        RECT 131.000 92.700 132.300 93.100 ;
        RECT 123.000 91.100 123.400 92.500 ;
        RECT 123.800 91.100 124.200 92.500 ;
        RECT 124.600 91.100 125.000 92.500 ;
        RECT 125.400 91.100 125.800 92.500 ;
        RECT 127.000 91.100 127.400 92.500 ;
        RECT 128.600 91.100 129.000 92.500 ;
        RECT 129.400 91.100 129.800 92.500 ;
        RECT 130.200 91.100 130.600 92.500 ;
        RECT 131.000 91.100 131.400 92.700 ;
        RECT 134.200 91.100 134.600 94.100 ;
        RECT 136.600 97.300 137.600 97.600 ;
        RECT 136.600 94.500 137.000 97.300 ;
        RECT 137.900 97.200 140.000 97.600 ;
        RECT 142.200 97.500 142.600 99.900 ;
        RECT 143.800 97.500 144.200 99.900 ;
        RECT 137.900 97.000 138.200 97.200 ;
        RECT 137.400 96.600 138.200 97.000 ;
        RECT 139.700 96.900 142.600 97.200 ;
        RECT 138.700 96.600 139.400 96.900 ;
        RECT 138.700 96.500 141.800 96.600 ;
        RECT 139.100 96.300 141.800 96.500 ;
        RECT 141.400 96.200 141.800 96.300 ;
        RECT 142.300 96.500 142.600 96.900 ;
        RECT 142.900 96.800 144.200 97.200 ;
        RECT 145.400 96.800 145.800 99.900 ;
        RECT 146.200 98.500 146.600 99.900 ;
        RECT 147.000 98.500 147.400 99.900 ;
        RECT 147.800 98.500 148.200 99.900 ;
        RECT 147.000 97.200 149.100 97.600 ;
        RECT 149.400 97.200 149.800 99.900 ;
        RECT 151.000 97.600 151.400 99.900 ;
        RECT 151.000 97.300 152.300 97.600 ;
        RECT 149.400 96.800 150.700 97.200 ;
        RECT 146.200 96.500 146.600 96.600 ;
        RECT 142.300 96.200 146.600 96.500 ;
        RECT 147.800 96.500 148.200 96.600 ;
        RECT 152.000 96.500 152.300 97.300 ;
        RECT 147.800 96.200 152.300 96.500 ;
        RECT 152.000 95.300 152.300 96.200 ;
        RECT 152.600 96.000 153.000 99.900 ;
        RECT 156.100 99.200 156.500 99.900 ;
        RECT 155.800 98.800 156.500 99.200 ;
        RECT 156.100 96.400 156.500 98.800 ;
        RECT 158.200 97.500 158.600 99.500 ;
        RECT 155.700 96.100 156.500 96.400 ;
        RECT 152.600 95.600 153.100 96.000 ;
        RECT 152.000 95.000 152.400 95.300 ;
        RECT 136.600 94.100 141.000 94.500 ;
        RECT 141.300 94.300 142.300 94.700 ;
        RECT 144.200 94.300 145.800 94.700 ;
        RECT 136.600 91.100 137.000 94.100 ;
        RECT 137.800 93.400 139.300 93.800 ;
        RECT 138.900 93.100 139.300 93.400 ;
        RECT 141.900 93.100 142.300 94.300 ;
        RECT 143.000 93.400 143.400 94.200 ;
        RECT 145.600 93.900 146.000 94.000 ;
        RECT 143.800 93.600 146.000 93.900 ;
        RECT 143.800 93.500 144.200 93.600 ;
        RECT 147.000 93.200 147.400 94.600 ;
        RECT 149.900 94.300 151.800 94.700 ;
        RECT 149.900 93.700 150.300 94.300 ;
        RECT 152.100 94.000 152.400 95.000 ;
        RECT 143.800 93.100 144.200 93.200 ;
        RECT 138.900 92.700 140.200 93.100 ;
        RECT 141.900 92.800 144.200 93.100 ;
        RECT 144.600 92.800 145.400 93.200 ;
        RECT 146.900 92.800 147.400 93.200 ;
        RECT 149.400 93.400 150.300 93.700 ;
        RECT 151.800 93.700 152.400 94.000 ;
        RECT 149.400 93.100 149.800 93.400 ;
        RECT 139.800 91.100 140.200 92.700 ;
        RECT 148.600 92.700 149.800 93.100 ;
        RECT 140.600 91.100 141.000 92.500 ;
        RECT 141.400 91.100 141.800 92.500 ;
        RECT 142.200 91.100 142.600 92.500 ;
        RECT 143.800 91.100 144.200 92.500 ;
        RECT 145.400 91.100 145.800 92.500 ;
        RECT 146.200 91.100 146.600 92.500 ;
        RECT 147.000 91.100 147.400 92.500 ;
        RECT 147.800 91.100 148.200 92.500 ;
        RECT 148.600 91.100 149.000 92.700 ;
        RECT 151.800 91.100 152.200 93.700 ;
        RECT 152.700 93.400 153.100 95.600 ;
        RECT 155.000 94.800 155.400 95.600 ;
        RECT 155.700 94.200 156.000 96.100 ;
        RECT 158.300 95.800 158.600 97.500 ;
        RECT 160.900 96.400 161.300 99.900 ;
        RECT 163.000 97.500 163.400 99.500 ;
        RECT 156.700 95.500 158.600 95.800 ;
        RECT 160.500 96.100 161.300 96.400 ;
        RECT 160.500 95.800 161.000 96.100 ;
        RECT 163.100 95.800 163.400 97.500 ;
        RECT 156.700 94.500 157.000 95.500 ;
        RECT 155.000 93.800 156.000 94.200 ;
        RECT 156.300 94.100 157.000 94.500 ;
        RECT 157.400 94.400 157.800 95.200 ;
        RECT 158.200 94.400 158.600 95.200 ;
        RECT 159.800 94.800 160.200 95.600 ;
        RECT 160.500 94.200 160.800 95.800 ;
        RECT 161.500 95.500 163.400 95.800 ;
        RECT 161.500 94.500 161.800 95.500 ;
        RECT 152.600 93.000 153.100 93.400 ;
        RECT 155.700 93.500 156.000 93.800 ;
        RECT 156.500 93.900 157.000 94.100 ;
        RECT 156.500 93.600 158.600 93.900 ;
        RECT 159.800 93.800 160.800 94.200 ;
        RECT 161.100 94.100 161.800 94.500 ;
        RECT 162.200 94.400 162.600 95.200 ;
        RECT 163.000 94.400 163.400 95.200 ;
        RECT 163.800 95.100 164.200 99.900 ;
        RECT 165.400 95.600 165.800 99.900 ;
        RECT 167.500 97.900 168.100 99.900 ;
        RECT 169.800 97.900 170.200 99.900 ;
        RECT 172.000 98.200 172.400 99.900 ;
        RECT 172.000 97.900 173.000 98.200 ;
        RECT 167.800 97.500 168.200 97.900 ;
        RECT 169.900 97.600 170.200 97.900 ;
        RECT 169.500 97.300 171.300 97.600 ;
        RECT 172.600 97.500 173.000 97.900 ;
        RECT 169.500 97.200 169.900 97.300 ;
        RECT 170.900 97.200 171.300 97.300 ;
        RECT 167.400 96.600 168.100 97.000 ;
        RECT 167.800 96.100 168.100 96.600 ;
        RECT 168.900 96.500 170.000 96.800 ;
        RECT 168.900 96.400 169.300 96.500 ;
        RECT 167.800 95.800 169.000 96.100 ;
        RECT 165.400 95.300 167.500 95.600 ;
        RECT 164.600 95.100 165.000 95.200 ;
        RECT 163.800 94.800 165.000 95.100 ;
        RECT 155.700 93.300 156.100 93.500 ;
        RECT 155.700 93.000 156.500 93.300 ;
        RECT 152.600 91.100 153.000 93.000 ;
        RECT 156.100 91.500 156.500 93.000 ;
        RECT 158.300 92.500 158.600 93.600 ;
        RECT 160.500 93.500 160.800 93.800 ;
        RECT 161.300 93.900 161.800 94.100 ;
        RECT 161.300 93.600 163.400 93.900 ;
        RECT 160.500 93.300 160.900 93.500 ;
        RECT 160.500 93.000 161.300 93.300 ;
        RECT 158.200 91.500 158.600 92.500 ;
        RECT 160.900 91.500 161.300 93.000 ;
        RECT 163.100 92.500 163.400 93.600 ;
        RECT 163.000 91.500 163.400 92.500 ;
        RECT 163.800 91.100 164.200 94.800 ;
        RECT 165.400 93.600 165.800 95.300 ;
        RECT 167.100 95.200 167.500 95.300 ;
        RECT 166.300 94.900 166.700 95.000 ;
        RECT 166.300 94.600 168.200 94.900 ;
        RECT 167.800 94.500 168.200 94.600 ;
        RECT 168.700 94.200 169.000 95.800 ;
        RECT 169.700 95.900 170.000 96.500 ;
        RECT 170.300 96.500 170.700 96.600 ;
        RECT 172.600 96.500 173.000 96.600 ;
        RECT 170.300 96.200 173.000 96.500 ;
        RECT 169.700 95.700 172.100 95.900 ;
        RECT 174.200 95.700 174.600 99.900 ;
        RECT 175.000 96.200 175.400 99.900 ;
        RECT 177.400 96.200 177.800 99.900 ;
        RECT 175.000 95.900 176.100 96.200 ;
        RECT 177.400 95.900 178.500 96.200 ;
        RECT 169.700 95.600 174.600 95.700 ;
        RECT 171.700 95.500 174.600 95.600 ;
        RECT 171.800 95.400 174.600 95.500 ;
        RECT 175.800 95.600 176.100 95.900 ;
        RECT 178.200 95.600 178.500 95.900 ;
        RECT 175.800 95.200 176.400 95.600 ;
        RECT 178.200 95.200 178.800 95.600 ;
        RECT 171.000 95.100 171.400 95.200 ;
        RECT 171.000 94.800 173.500 95.100 ;
        RECT 173.100 94.700 173.500 94.800 ;
        RECT 175.000 94.400 175.400 95.200 ;
        RECT 172.300 94.200 172.700 94.300 ;
        RECT 168.700 93.900 174.200 94.200 ;
        RECT 168.900 93.800 169.300 93.900 ;
        RECT 165.400 93.300 167.300 93.600 ;
        RECT 164.600 93.100 165.000 93.200 ;
        RECT 165.400 93.100 165.800 93.300 ;
        RECT 166.900 93.200 167.300 93.300 ;
        RECT 164.600 92.800 165.800 93.100 ;
        RECT 171.800 92.800 172.100 93.900 ;
        RECT 173.400 93.800 174.200 93.900 ;
        RECT 175.800 93.700 176.100 95.200 ;
        RECT 177.400 94.400 177.800 95.200 ;
        RECT 178.200 93.700 178.500 95.200 ;
        RECT 164.600 92.400 165.000 92.800 ;
        RECT 165.400 91.100 165.800 92.800 ;
        RECT 170.900 92.700 171.300 92.800 ;
        RECT 167.800 92.100 168.200 92.500 ;
        RECT 169.900 92.400 171.300 92.700 ;
        RECT 171.800 92.400 172.200 92.800 ;
        RECT 169.900 92.100 170.200 92.400 ;
        RECT 172.600 92.100 173.000 92.500 ;
        RECT 167.500 91.800 168.200 92.100 ;
        RECT 167.500 91.100 168.100 91.800 ;
        RECT 169.800 91.100 170.200 92.100 ;
        RECT 172.000 91.800 173.000 92.100 ;
        RECT 172.000 91.100 172.400 91.800 ;
        RECT 174.200 91.100 174.600 93.500 ;
        RECT 175.000 93.400 176.100 93.700 ;
        RECT 177.400 93.400 178.500 93.700 ;
        RECT 175.000 91.100 175.400 93.400 ;
        RECT 177.400 91.100 177.800 93.400 ;
        RECT 0.600 87.500 1.000 89.900 ;
        RECT 2.800 89.200 3.200 89.900 ;
        RECT 2.200 88.900 3.200 89.200 ;
        RECT 5.000 88.900 5.400 89.900 ;
        RECT 7.100 89.200 7.700 89.900 ;
        RECT 7.000 88.900 7.700 89.200 ;
        RECT 2.200 88.500 2.600 88.900 ;
        RECT 5.000 88.600 5.300 88.900 ;
        RECT 3.000 87.800 3.400 88.600 ;
        RECT 3.900 88.300 5.300 88.600 ;
        RECT 7.000 88.500 7.400 88.900 ;
        RECT 3.900 88.200 4.300 88.300 ;
        RECT 1.000 87.100 1.800 87.200 ;
        RECT 3.100 87.100 3.400 87.800 ;
        RECT 7.900 87.700 8.300 87.800 ;
        RECT 9.400 87.700 9.800 89.900 ;
        RECT 10.300 88.200 10.700 88.600 ;
        RECT 10.200 87.800 10.600 88.200 ;
        RECT 11.000 87.900 11.400 89.900 ;
        RECT 14.200 88.900 14.600 89.900 ;
        RECT 7.900 87.400 9.800 87.700 ;
        RECT 5.900 87.100 6.300 87.200 ;
        RECT 1.000 86.800 6.500 87.100 ;
        RECT 2.500 86.700 2.900 86.800 ;
        RECT 1.700 86.200 2.100 86.300 ;
        RECT 6.200 86.200 6.500 86.800 ;
        RECT 7.000 86.400 7.400 86.500 ;
        RECT 1.700 85.900 4.200 86.200 ;
        RECT 3.800 85.800 4.200 85.900 ;
        RECT 6.200 85.800 6.600 86.200 ;
        RECT 7.000 86.100 8.900 86.400 ;
        RECT 8.500 86.000 8.900 86.100 ;
        RECT 0.600 85.500 3.400 85.600 ;
        RECT 0.600 85.400 3.500 85.500 ;
        RECT 0.600 85.300 5.500 85.400 ;
        RECT 0.600 81.100 1.000 85.300 ;
        RECT 3.100 85.100 5.500 85.300 ;
        RECT 2.200 84.500 4.900 84.800 ;
        RECT 2.200 84.400 2.600 84.500 ;
        RECT 4.500 84.400 4.900 84.500 ;
        RECT 5.200 84.500 5.500 85.100 ;
        RECT 6.200 85.200 6.500 85.800 ;
        RECT 7.700 85.700 8.100 85.800 ;
        RECT 9.400 85.700 9.800 87.400 ;
        RECT 10.200 86.800 10.600 87.200 ;
        RECT 10.200 86.200 10.500 86.800 ;
        RECT 10.200 86.100 10.600 86.200 ;
        RECT 11.100 86.100 11.400 87.900 ;
        RECT 13.400 88.100 13.800 88.200 ;
        RECT 14.200 88.100 14.500 88.900 ;
        RECT 13.400 87.800 14.500 88.100 ;
        RECT 14.200 87.200 14.500 87.800 ;
        RECT 15.000 87.800 15.400 88.600 ;
        RECT 17.100 88.200 17.500 89.900 ;
        RECT 18.500 89.200 18.900 89.900 ;
        RECT 18.200 88.800 18.900 89.200 ;
        RECT 18.500 88.400 18.900 88.800 ;
        RECT 16.600 87.900 17.500 88.200 ;
        RECT 18.200 87.900 18.900 88.400 ;
        RECT 20.600 87.900 21.000 89.900 ;
        RECT 22.700 88.200 23.100 89.900 ;
        RECT 22.200 87.900 23.100 88.200 ;
        RECT 24.400 89.100 24.800 89.900 ;
        RECT 24.400 88.800 25.700 89.100 ;
        RECT 11.800 87.100 12.200 87.200 ;
        RECT 11.800 86.800 13.700 87.100 ;
        RECT 11.800 86.400 12.200 86.800 ;
        RECT 13.400 86.200 13.700 86.800 ;
        RECT 14.200 86.800 14.600 87.200 ;
        RECT 15.000 87.100 15.300 87.800 ;
        RECT 15.800 87.100 16.200 87.600 ;
        RECT 15.000 86.800 16.200 87.100 ;
        RECT 12.600 86.100 13.000 86.200 ;
        RECT 10.200 85.800 11.400 86.100 ;
        RECT 12.200 85.800 13.000 86.100 ;
        RECT 7.700 85.400 9.800 85.700 ;
        RECT 6.200 84.900 7.400 85.200 ;
        RECT 5.900 84.500 6.300 84.600 ;
        RECT 5.200 84.200 6.300 84.500 ;
        RECT 7.100 84.400 7.400 84.900 ;
        RECT 7.100 84.000 7.800 84.400 ;
        RECT 3.900 83.700 4.300 83.800 ;
        RECT 5.300 83.700 5.700 83.800 ;
        RECT 2.200 83.100 2.600 83.500 ;
        RECT 3.900 83.400 5.700 83.700 ;
        RECT 5.000 83.100 5.300 83.400 ;
        RECT 7.000 83.100 7.400 83.500 ;
        RECT 2.200 82.800 3.200 83.100 ;
        RECT 2.800 81.100 3.200 82.800 ;
        RECT 5.000 81.100 5.400 83.100 ;
        RECT 7.100 81.100 7.700 83.100 ;
        RECT 9.400 81.100 9.800 85.400 ;
        RECT 10.300 85.100 10.600 85.800 ;
        RECT 12.200 85.600 12.600 85.800 ;
        RECT 13.400 85.400 13.800 86.200 ;
        RECT 14.200 85.100 14.500 86.800 ;
        RECT 16.600 86.100 17.000 87.900 ;
        RECT 17.400 86.800 17.800 87.200 ;
        RECT 17.400 86.100 17.700 86.800 ;
        RECT 16.600 85.800 17.700 86.100 ;
        RECT 18.200 86.200 18.500 87.900 ;
        RECT 20.600 87.800 20.900 87.900 ;
        RECT 20.000 87.600 20.900 87.800 ;
        RECT 18.800 87.500 20.900 87.600 ;
        RECT 18.800 87.300 20.300 87.500 ;
        RECT 18.800 87.200 19.200 87.300 ;
        RECT 18.200 85.800 18.600 86.200 ;
        RECT 10.200 81.100 10.600 85.100 ;
        RECT 11.000 84.800 13.000 85.100 ;
        RECT 11.000 81.100 11.400 84.800 ;
        RECT 12.600 81.100 13.000 84.800 ;
        RECT 13.700 84.700 14.600 85.100 ;
        RECT 13.700 81.100 14.100 84.700 ;
        RECT 16.600 81.100 17.000 85.800 ;
        RECT 17.400 84.400 17.800 85.200 ;
        RECT 18.200 85.100 18.500 85.800 ;
        RECT 18.900 85.500 19.200 87.200 ;
        RECT 19.600 86.900 20.000 87.000 ;
        RECT 19.600 86.600 20.100 86.900 ;
        RECT 19.800 86.200 20.100 86.600 ;
        RECT 20.600 86.400 21.000 87.200 ;
        RECT 21.400 86.800 21.800 87.600 ;
        RECT 19.800 85.800 20.200 86.200 ;
        RECT 18.900 85.200 20.100 85.500 ;
        RECT 18.200 81.100 18.600 85.100 ;
        RECT 19.800 83.100 20.100 85.200 ;
        RECT 19.800 81.100 20.200 83.100 ;
        RECT 22.200 81.100 22.600 87.900 ;
        RECT 24.400 87.100 24.800 88.800 ;
        RECT 25.400 88.200 25.700 88.800 ;
        RECT 27.300 88.200 27.700 89.900 ;
        RECT 31.000 89.200 31.400 89.900 ;
        RECT 31.000 88.900 31.500 89.200 ;
        RECT 31.200 88.800 31.500 88.900 ;
        RECT 32.600 88.900 33.000 89.900 ;
        RECT 32.600 88.800 33.200 88.900 ;
        RECT 31.200 88.500 33.200 88.800 ;
        RECT 25.400 87.800 25.800 88.200 ;
        RECT 27.300 87.900 28.200 88.200 ;
        RECT 23.900 86.900 24.800 87.100 ;
        RECT 23.900 86.800 24.700 86.900 ;
        RECT 23.900 85.200 24.200 86.800 ;
        RECT 25.000 85.800 25.800 86.200 ;
        RECT 23.000 84.400 23.400 85.200 ;
        RECT 23.800 84.800 24.200 85.200 ;
        RECT 26.200 84.800 26.600 85.600 ;
        RECT 23.900 83.500 24.200 84.800 ;
        RECT 24.600 83.800 25.000 84.600 ;
        RECT 27.000 84.400 27.400 85.200 ;
        RECT 23.900 83.200 25.700 83.500 ;
        RECT 23.900 83.100 24.200 83.200 ;
        RECT 23.800 81.100 24.200 83.100 ;
        RECT 25.400 83.100 25.700 83.200 ;
        RECT 25.400 81.100 25.800 83.100 ;
        RECT 27.800 81.100 28.200 87.900 ;
        RECT 30.200 87.800 31.100 88.200 ;
        RECT 28.600 87.100 29.000 87.600 ;
        RECT 29.400 87.100 29.800 87.200 ;
        RECT 28.600 86.800 29.800 87.100 ;
        RECT 31.000 86.800 31.800 87.200 ;
        RECT 28.600 86.100 29.000 86.200 ;
        RECT 31.000 86.100 31.300 86.800 ;
        RECT 28.600 85.800 31.300 86.100 ;
        RECT 31.800 85.800 32.600 86.200 ;
        RECT 32.900 85.200 33.200 88.500 ;
        RECT 37.600 87.100 38.000 89.900 ;
        RECT 41.900 87.900 42.700 89.900 ;
        RECT 45.900 89.200 46.300 89.900 ;
        RECT 45.400 88.800 46.300 89.200 ;
        RECT 45.900 88.200 46.300 88.800 ;
        RECT 45.400 87.900 46.300 88.200 ;
        RECT 39.000 87.100 39.400 87.200 ;
        RECT 41.400 87.100 41.800 87.200 ;
        RECT 37.600 86.900 38.500 87.100 ;
        RECT 37.700 86.800 38.500 86.900 ;
        RECT 39.000 86.800 41.800 87.100 ;
        RECT 34.200 85.600 36.100 85.900 ;
        RECT 36.600 85.800 37.800 86.200 ;
        RECT 34.200 85.500 34.600 85.600 ;
        RECT 32.900 85.100 34.600 85.200 ;
        RECT 35.000 85.100 35.400 85.200 ;
        RECT 32.900 84.900 35.400 85.100 ;
        RECT 34.200 84.800 35.400 84.900 ;
        RECT 35.800 84.800 36.200 85.600 ;
        RECT 38.200 85.200 38.500 86.800 ;
        RECT 41.500 86.600 41.800 86.800 ;
        RECT 41.500 86.200 41.900 86.600 ;
        RECT 42.200 86.200 42.500 87.900 ;
        RECT 43.000 86.400 43.400 87.200 ;
        RECT 44.600 86.800 45.000 87.600 ;
        RECT 40.600 85.400 41.000 86.200 ;
        RECT 42.200 85.800 42.600 86.200 ;
        RECT 43.800 86.100 44.200 86.200 ;
        RECT 43.400 85.800 44.200 86.100 ;
        RECT 42.200 85.700 42.500 85.800 ;
        RECT 41.500 85.400 42.500 85.700 ;
        RECT 43.400 85.600 43.800 85.800 ;
        RECT 38.200 84.800 38.600 85.200 ;
        RECT 41.500 85.100 41.800 85.400 ;
        RECT 29.500 84.400 31.300 84.700 ;
        RECT 29.500 84.100 29.800 84.400 ;
        RECT 29.400 81.100 29.800 84.100 ;
        RECT 31.000 84.100 31.300 84.400 ;
        RECT 31.900 84.500 33.700 84.600 ;
        RECT 34.200 84.500 34.500 84.800 ;
        RECT 31.900 84.300 33.800 84.500 ;
        RECT 31.900 84.100 32.200 84.300 ;
        RECT 31.000 81.400 31.400 84.100 ;
        RECT 31.800 81.700 32.200 84.100 ;
        RECT 32.600 81.400 33.000 84.000 ;
        RECT 33.400 81.500 33.800 84.300 ;
        RECT 34.200 81.700 34.600 84.500 ;
        RECT 31.000 81.100 33.000 81.400 ;
        RECT 33.500 81.400 33.800 81.500 ;
        RECT 35.000 81.500 35.400 84.500 ;
        RECT 36.600 84.100 37.000 84.200 ;
        RECT 37.400 84.100 37.800 84.600 ;
        RECT 36.600 83.800 37.800 84.100 ;
        RECT 38.200 83.500 38.500 84.800 ;
        RECT 36.700 83.200 38.500 83.500 ;
        RECT 36.700 83.100 37.000 83.200 ;
        RECT 35.000 81.400 35.300 81.500 ;
        RECT 33.500 81.100 35.300 81.400 ;
        RECT 36.600 81.100 37.000 83.100 ;
        RECT 38.200 83.100 38.500 83.200 ;
        RECT 38.200 82.100 38.600 83.100 ;
        RECT 39.000 82.100 39.400 82.200 ;
        RECT 38.200 81.800 39.400 82.100 ;
        RECT 38.200 81.100 38.600 81.800 ;
        RECT 40.600 81.400 41.000 85.100 ;
        RECT 41.400 81.700 41.800 85.100 ;
        RECT 42.200 84.800 44.200 85.100 ;
        RECT 42.200 81.400 42.600 84.800 ;
        RECT 40.600 81.100 42.600 81.400 ;
        RECT 43.800 81.100 44.200 84.800 ;
        RECT 45.400 81.100 45.800 87.900 ;
        RECT 47.000 87.700 47.400 89.900 ;
        RECT 49.100 89.200 49.700 89.900 ;
        RECT 49.100 88.900 49.800 89.200 ;
        RECT 51.400 88.900 51.800 89.900 ;
        RECT 53.600 89.200 54.000 89.900 ;
        RECT 53.600 88.900 54.600 89.200 ;
        RECT 49.400 88.500 49.800 88.900 ;
        RECT 51.500 88.600 51.800 88.900 ;
        RECT 51.500 88.300 52.900 88.600 ;
        RECT 52.500 88.200 52.900 88.300 ;
        RECT 53.400 88.200 53.800 88.600 ;
        RECT 54.200 88.500 54.600 88.900 ;
        RECT 48.500 87.700 48.900 87.800 ;
        RECT 47.000 87.400 48.900 87.700 ;
        RECT 47.000 85.700 47.400 87.400 ;
        RECT 50.500 87.100 50.900 87.200 ;
        RECT 53.400 87.100 53.700 88.200 ;
        RECT 55.800 87.500 56.200 89.900 ;
        RECT 58.200 87.900 58.600 89.900 ;
        RECT 60.600 88.900 61.000 89.900 ;
        RECT 58.900 88.200 59.300 88.600 ;
        RECT 55.000 87.100 55.800 87.200 ;
        RECT 50.300 86.800 55.800 87.100 ;
        RECT 49.400 86.400 49.800 86.500 ;
        RECT 47.900 86.100 49.800 86.400 ;
        RECT 47.900 86.000 48.300 86.100 ;
        RECT 48.700 85.700 49.100 85.800 ;
        RECT 47.000 85.400 49.100 85.700 ;
        RECT 46.200 84.400 46.600 85.200 ;
        RECT 47.000 81.100 47.400 85.400 ;
        RECT 50.300 85.200 50.600 86.800 ;
        RECT 53.900 86.700 54.300 86.800 ;
        RECT 57.400 86.400 57.800 87.200 ;
        RECT 53.400 86.200 53.800 86.300 ;
        RECT 54.700 86.200 55.100 86.300 ;
        RECT 52.600 85.900 55.100 86.200 ;
        RECT 56.600 86.100 57.000 86.200 ;
        RECT 58.200 86.100 58.500 87.900 ;
        RECT 59.000 87.800 59.400 88.200 ;
        RECT 59.800 87.800 60.200 88.600 ;
        RECT 59.000 87.100 59.300 87.800 ;
        RECT 60.700 87.200 61.000 88.900 ;
        RECT 63.500 88.200 63.900 89.900 ;
        RECT 65.200 89.200 65.600 89.900 ;
        RECT 64.600 88.800 65.600 89.200 ;
        RECT 63.000 87.900 63.900 88.200 ;
        RECT 60.600 87.100 61.000 87.200 ;
        RECT 59.000 86.800 61.000 87.100 ;
        RECT 62.200 86.800 62.600 87.600 ;
        RECT 59.000 86.100 59.400 86.200 ;
        RECT 52.600 85.800 53.000 85.900 ;
        RECT 56.600 85.800 57.400 86.100 ;
        RECT 58.200 85.800 59.400 86.100 ;
        RECT 57.000 85.600 57.400 85.800 ;
        RECT 53.400 85.500 56.200 85.600 ;
        RECT 53.300 85.400 56.200 85.500 ;
        RECT 49.400 84.900 50.600 85.200 ;
        RECT 51.300 85.300 56.200 85.400 ;
        RECT 51.300 85.100 53.700 85.300 ;
        RECT 49.400 84.400 49.700 84.900 ;
        RECT 49.000 84.000 49.700 84.400 ;
        RECT 50.500 84.500 50.900 84.600 ;
        RECT 51.300 84.500 51.600 85.100 ;
        RECT 50.500 84.200 51.600 84.500 ;
        RECT 51.900 84.500 54.600 84.800 ;
        RECT 51.900 84.400 52.300 84.500 ;
        RECT 54.200 84.400 54.600 84.500 ;
        RECT 51.100 83.700 51.500 83.800 ;
        RECT 52.500 83.700 52.900 83.800 ;
        RECT 49.400 83.100 49.800 83.500 ;
        RECT 51.100 83.400 52.900 83.700 ;
        RECT 51.500 83.100 51.800 83.400 ;
        RECT 54.200 83.100 54.600 83.500 ;
        RECT 49.100 81.100 49.700 83.100 ;
        RECT 51.400 81.100 51.800 83.100 ;
        RECT 53.600 82.800 54.600 83.100 ;
        RECT 53.600 81.100 54.000 82.800 ;
        RECT 55.800 81.100 56.200 85.300 ;
        RECT 59.000 85.100 59.300 85.800 ;
        RECT 60.700 85.100 61.000 86.800 ;
        RECT 61.400 85.400 61.800 86.200 ;
        RECT 56.600 84.800 58.600 85.100 ;
        RECT 56.600 81.100 57.000 84.800 ;
        RECT 58.200 81.100 58.600 84.800 ;
        RECT 59.000 81.100 59.400 85.100 ;
        RECT 60.600 84.700 61.500 85.100 ;
        RECT 61.100 81.100 61.500 84.700 ;
        RECT 63.000 81.100 63.400 87.900 ;
        RECT 65.200 87.100 65.600 88.800 ;
        RECT 69.100 88.200 69.500 89.900 ;
        RECT 71.000 88.900 71.400 89.900 ;
        RECT 68.600 87.800 69.700 88.200 ;
        RECT 70.200 87.800 70.600 88.600 ;
        RECT 71.100 88.100 71.400 88.900 ;
        RECT 72.700 88.200 73.100 88.600 ;
        RECT 72.600 88.100 73.000 88.200 ;
        RECT 71.000 87.800 73.000 88.100 ;
        RECT 73.400 87.900 73.800 89.900 ;
        RECT 64.700 86.900 65.600 87.100 ;
        RECT 64.700 86.800 65.500 86.900 ;
        RECT 67.800 86.800 68.200 87.600 ;
        RECT 64.700 85.200 65.000 86.800 ;
        RECT 65.800 85.800 66.600 86.200 ;
        RECT 67.000 85.800 68.100 86.100 ;
        RECT 63.800 84.400 64.200 85.200 ;
        RECT 64.600 84.800 65.000 85.200 ;
        RECT 67.000 84.800 67.400 85.800 ;
        RECT 67.800 85.200 68.100 85.800 ;
        RECT 67.800 84.800 68.200 85.200 ;
        RECT 64.700 83.500 65.000 84.800 ;
        RECT 65.400 83.800 65.800 84.600 ;
        RECT 64.700 83.200 66.500 83.500 ;
        RECT 64.700 83.100 65.000 83.200 ;
        RECT 64.600 81.100 65.000 83.100 ;
        RECT 66.200 83.100 66.500 83.200 ;
        RECT 66.200 81.100 66.600 83.100 ;
        RECT 68.600 81.100 69.000 87.800 ;
        RECT 69.400 87.200 69.700 87.800 ;
        RECT 71.100 87.200 71.400 87.800 ;
        RECT 69.400 86.800 69.800 87.200 ;
        RECT 71.000 86.800 71.400 87.200 ;
        RECT 69.400 84.400 69.800 85.200 ;
        RECT 71.100 85.100 71.400 86.800 ;
        RECT 71.800 85.400 72.200 86.200 ;
        RECT 72.600 86.100 73.000 86.200 ;
        RECT 73.500 86.100 73.800 87.900 ;
        RECT 75.800 88.500 76.200 89.500 ;
        RECT 75.800 87.400 76.100 88.500 ;
        RECT 77.900 88.000 78.300 89.500 ;
        RECT 80.900 88.200 81.300 89.900 ;
        RECT 84.300 89.200 84.700 89.900 ;
        RECT 84.300 88.800 85.000 89.200 ;
        RECT 84.300 88.200 84.700 88.800 ;
        RECT 77.900 87.700 78.700 88.000 ;
        RECT 80.900 87.900 81.800 88.200 ;
        RECT 78.300 87.500 78.700 87.700 ;
        RECT 74.200 86.400 74.600 87.200 ;
        RECT 75.800 87.100 77.900 87.400 ;
        RECT 77.400 86.900 77.900 87.100 ;
        RECT 78.400 87.200 78.700 87.500 ;
        RECT 75.000 86.100 75.400 86.200 ;
        RECT 72.600 85.800 73.800 86.100 ;
        RECT 74.600 85.800 75.400 86.100 ;
        RECT 75.800 85.800 76.200 86.600 ;
        RECT 76.600 85.800 77.000 86.600 ;
        RECT 77.400 86.500 78.100 86.900 ;
        RECT 78.400 86.800 79.400 87.200 ;
        RECT 79.800 87.100 80.200 87.200 ;
        RECT 81.400 87.100 81.800 87.900 ;
        RECT 83.800 87.900 84.700 88.200 ;
        RECT 79.800 86.800 81.800 87.100 ;
        RECT 82.200 86.800 82.600 87.600 ;
        RECT 83.000 86.800 83.400 87.600 ;
        RECT 72.700 85.100 73.000 85.800 ;
        RECT 74.600 85.600 75.000 85.800 ;
        RECT 77.400 85.500 77.700 86.500 ;
        RECT 75.800 85.200 77.700 85.500 ;
        RECT 71.000 84.700 71.900 85.100 ;
        RECT 71.500 81.100 71.900 84.700 ;
        RECT 72.600 81.100 73.000 85.100 ;
        RECT 73.400 84.800 75.400 85.100 ;
        RECT 73.400 81.100 73.800 84.800 ;
        RECT 75.000 81.100 75.400 84.800 ;
        RECT 75.800 83.500 76.100 85.200 ;
        RECT 78.400 84.900 78.700 86.800 ;
        RECT 79.000 85.400 79.400 86.200 ;
        RECT 77.900 84.600 78.700 84.900 ;
        RECT 75.800 81.500 76.200 83.500 ;
        RECT 77.900 82.200 78.300 84.600 ;
        RECT 80.600 84.400 81.000 85.200 ;
        RECT 77.900 81.800 78.600 82.200 ;
        RECT 77.900 81.100 78.300 81.800 ;
        RECT 81.400 81.100 81.800 86.800 ;
        RECT 83.800 81.100 84.200 87.900 ;
        RECT 85.400 87.800 85.800 88.600 ;
        RECT 86.200 86.100 86.600 89.900 ;
        RECT 90.500 89.200 90.900 89.500 ;
        RECT 90.500 88.800 91.400 89.200 ;
        RECT 90.500 88.000 90.900 88.800 ;
        RECT 92.600 88.500 93.000 89.500 ;
        RECT 94.200 88.900 94.600 89.900 ;
        RECT 90.100 87.700 90.900 88.000 ;
        RECT 90.100 87.500 90.500 87.700 ;
        RECT 90.100 87.200 90.400 87.500 ;
        RECT 92.700 87.400 93.000 88.500 ;
        RECT 93.400 87.800 93.800 88.600 ;
        RECT 94.300 88.100 94.600 88.900 ;
        RECT 95.900 88.200 96.300 88.600 ;
        RECT 95.800 88.100 96.200 88.200 ;
        RECT 94.200 87.800 96.200 88.100 ;
        RECT 96.600 87.900 97.000 89.900 ;
        RECT 100.900 88.200 101.300 89.500 ;
        RECT 103.000 88.500 103.400 89.500 ;
        RECT 100.900 88.000 101.800 88.200 ;
        RECT 89.400 86.800 90.400 87.200 ;
        RECT 90.900 87.100 93.000 87.400 ;
        RECT 94.300 87.200 94.600 87.800 ;
        RECT 90.900 86.900 91.400 87.100 ;
        RECT 89.400 86.100 89.800 86.200 ;
        RECT 86.200 85.800 89.800 86.100 ;
        RECT 84.600 84.400 85.000 85.200 ;
        RECT 86.200 81.100 86.600 85.800 ;
        RECT 89.400 85.400 89.800 85.800 ;
        RECT 90.100 84.900 90.400 86.800 ;
        RECT 90.700 86.500 91.400 86.900 ;
        RECT 94.200 86.800 94.600 87.200 ;
        RECT 91.100 85.500 91.400 86.500 ;
        RECT 91.800 85.800 92.200 86.600 ;
        RECT 92.600 86.100 93.000 86.600 ;
        RECT 93.400 86.100 93.800 86.200 ;
        RECT 92.600 85.800 93.800 86.100 ;
        RECT 91.100 85.200 93.000 85.500 ;
        RECT 90.100 84.600 90.900 84.900 ;
        RECT 90.500 81.100 90.900 84.600 ;
        RECT 92.700 83.500 93.000 85.200 ;
        RECT 94.300 85.100 94.600 86.800 ;
        RECT 95.000 85.400 95.400 86.200 ;
        RECT 95.800 86.100 96.200 86.200 ;
        RECT 96.700 86.100 97.000 87.900 ;
        RECT 100.500 87.800 101.800 88.000 ;
        RECT 100.500 87.700 101.300 87.800 ;
        RECT 100.500 87.500 100.900 87.700 ;
        RECT 100.500 87.200 100.800 87.500 ;
        RECT 103.100 87.400 103.400 88.500 ;
        RECT 103.800 87.500 104.200 89.900 ;
        RECT 106.000 89.200 106.400 89.900 ;
        RECT 105.400 88.900 106.400 89.200 ;
        RECT 108.200 88.900 108.600 89.900 ;
        RECT 110.300 89.200 110.900 89.900 ;
        RECT 110.200 88.900 110.900 89.200 ;
        RECT 105.400 88.500 105.800 88.900 ;
        RECT 108.200 88.600 108.500 88.900 ;
        RECT 106.200 87.800 106.600 88.600 ;
        RECT 107.100 88.300 108.500 88.600 ;
        RECT 110.200 88.500 110.600 88.900 ;
        RECT 107.100 88.200 107.500 88.300 ;
        RECT 112.600 88.100 113.000 89.900 ;
        RECT 113.400 88.100 113.800 88.600 ;
        RECT 112.600 87.800 113.800 88.100 ;
        RECT 97.400 87.100 97.800 87.200 ;
        RECT 99.000 87.100 99.400 87.200 ;
        RECT 97.400 86.800 99.400 87.100 ;
        RECT 99.800 86.800 100.800 87.200 ;
        RECT 101.300 87.100 103.400 87.400 ;
        RECT 104.200 87.100 105.000 87.200 ;
        RECT 106.300 87.100 106.600 87.800 ;
        RECT 111.100 87.700 111.500 87.800 ;
        RECT 112.600 87.700 113.000 87.800 ;
        RECT 111.100 87.400 113.000 87.700 ;
        RECT 109.100 87.100 109.500 87.200 ;
        RECT 101.300 86.900 101.800 87.100 ;
        RECT 97.400 86.400 97.800 86.800 ;
        RECT 98.200 86.100 98.600 86.200 ;
        RECT 95.800 85.800 97.000 86.100 ;
        RECT 97.800 85.800 98.600 86.100 ;
        RECT 95.900 85.100 96.200 85.800 ;
        RECT 97.800 85.600 98.200 85.800 ;
        RECT 99.800 85.400 100.200 86.200 ;
        RECT 94.200 84.700 95.100 85.100 ;
        RECT 92.600 81.500 93.000 83.500 ;
        RECT 94.700 81.100 95.100 84.700 ;
        RECT 95.800 81.100 96.200 85.100 ;
        RECT 96.600 84.800 98.600 85.100 ;
        RECT 96.600 81.100 97.000 84.800 ;
        RECT 98.200 81.100 98.600 84.800 ;
        RECT 100.500 84.900 100.800 86.800 ;
        RECT 101.100 86.500 101.800 86.900 ;
        RECT 104.200 86.800 109.700 87.100 ;
        RECT 105.700 86.700 106.100 86.800 ;
        RECT 101.500 85.500 101.800 86.500 ;
        RECT 102.200 85.800 102.600 86.600 ;
        RECT 103.000 85.800 103.400 86.600 ;
        RECT 104.900 86.200 105.300 86.300 ;
        RECT 106.200 86.200 106.600 86.300 ;
        RECT 104.900 85.900 107.400 86.200 ;
        RECT 107.000 85.800 107.400 85.900 ;
        RECT 103.800 85.500 106.600 85.600 ;
        RECT 101.500 85.200 103.400 85.500 ;
        RECT 100.500 84.600 101.300 84.900 ;
        RECT 100.900 81.100 101.300 84.600 ;
        RECT 103.100 83.500 103.400 85.200 ;
        RECT 103.000 81.500 103.400 83.500 ;
        RECT 103.800 85.400 106.700 85.500 ;
        RECT 103.800 85.300 108.700 85.400 ;
        RECT 103.800 81.100 104.200 85.300 ;
        RECT 106.300 85.100 108.700 85.300 ;
        RECT 105.400 84.500 108.100 84.800 ;
        RECT 105.400 84.400 105.800 84.500 ;
        RECT 107.700 84.400 108.100 84.500 ;
        RECT 108.400 84.500 108.700 85.100 ;
        RECT 109.400 85.200 109.700 86.800 ;
        RECT 110.200 86.400 110.600 86.500 ;
        RECT 110.200 86.100 112.100 86.400 ;
        RECT 111.700 86.000 112.100 86.100 ;
        RECT 110.900 85.700 111.300 85.800 ;
        RECT 112.600 85.700 113.000 87.400 ;
        RECT 110.900 85.400 113.000 85.700 ;
        RECT 109.400 84.900 110.600 85.200 ;
        RECT 109.100 84.500 109.500 84.600 ;
        RECT 108.400 84.200 109.500 84.500 ;
        RECT 110.300 84.400 110.600 84.900 ;
        RECT 110.300 84.000 111.000 84.400 ;
        RECT 107.100 83.700 107.500 83.800 ;
        RECT 108.500 83.700 108.900 83.800 ;
        RECT 105.400 83.100 105.800 83.500 ;
        RECT 107.100 83.400 108.900 83.700 ;
        RECT 108.200 83.100 108.500 83.400 ;
        RECT 110.200 83.100 110.600 83.500 ;
        RECT 105.400 82.800 106.400 83.100 ;
        RECT 106.000 81.100 106.400 82.800 ;
        RECT 108.200 81.100 108.600 83.100 ;
        RECT 110.300 81.100 110.900 83.100 ;
        RECT 112.600 81.100 113.000 85.400 ;
        RECT 114.200 81.100 114.600 89.900 ;
        RECT 115.100 88.200 115.500 88.600 ;
        RECT 115.000 87.800 115.400 88.200 ;
        RECT 115.800 87.900 116.200 89.900 ;
        RECT 120.100 89.200 120.500 89.500 ;
        RECT 120.100 88.800 121.000 89.200 ;
        RECT 120.100 88.000 120.500 88.800 ;
        RECT 122.200 88.500 122.600 89.500 ;
        RECT 115.000 86.100 115.400 86.200 ;
        RECT 115.900 86.100 116.200 87.900 ;
        RECT 119.700 87.700 120.500 88.000 ;
        RECT 119.700 87.500 120.100 87.700 ;
        RECT 119.700 87.200 120.000 87.500 ;
        RECT 122.300 87.400 122.600 88.500 ;
        RECT 116.600 86.400 117.000 87.200 ;
        RECT 119.000 86.800 120.000 87.200 ;
        RECT 120.500 87.100 122.600 87.400 ;
        RECT 120.500 86.900 121.000 87.100 ;
        RECT 117.400 86.100 117.800 86.200 ;
        RECT 115.000 85.800 116.200 86.100 ;
        RECT 117.000 85.800 117.800 86.100 ;
        RECT 115.100 85.100 115.400 85.800 ;
        RECT 117.000 85.600 117.400 85.800 ;
        RECT 119.000 85.400 119.400 86.200 ;
        RECT 115.000 81.100 115.400 85.100 ;
        RECT 115.800 84.800 117.800 85.100 ;
        RECT 115.800 81.100 116.200 84.800 ;
        RECT 117.400 81.100 117.800 84.800 ;
        RECT 119.700 84.900 120.000 86.800 ;
        RECT 120.300 86.500 121.000 86.900 ;
        RECT 120.700 85.500 121.000 86.500 ;
        RECT 121.400 85.800 121.800 86.600 ;
        RECT 122.200 85.800 122.600 86.600 ;
        RECT 120.700 85.200 122.600 85.500 ;
        RECT 119.700 84.600 120.500 84.900 ;
        RECT 120.100 81.100 120.500 84.600 ;
        RECT 122.300 83.500 122.600 85.200 ;
        RECT 122.200 81.500 122.600 83.500 ;
        RECT 123.000 85.100 123.400 89.900 ;
        RECT 123.800 87.800 124.200 88.600 ;
        RECT 124.600 87.500 125.000 89.900 ;
        RECT 126.800 89.200 127.200 89.900 ;
        RECT 126.200 88.900 127.200 89.200 ;
        RECT 129.000 88.900 129.400 89.900 ;
        RECT 131.100 89.200 131.700 89.900 ;
        RECT 131.000 88.900 131.700 89.200 ;
        RECT 126.200 88.500 126.600 88.900 ;
        RECT 129.000 88.600 129.300 88.900 ;
        RECT 127.000 87.800 127.400 88.600 ;
        RECT 127.900 88.300 129.300 88.600 ;
        RECT 131.000 88.500 131.400 88.900 ;
        RECT 127.900 88.200 128.300 88.300 ;
        RECT 125.000 87.100 125.800 87.200 ;
        RECT 127.100 87.100 127.400 87.800 ;
        RECT 131.900 87.700 132.300 87.800 ;
        RECT 133.400 87.700 133.800 89.900 ;
        RECT 131.900 87.400 133.800 87.700 ;
        RECT 129.900 87.100 130.300 87.200 ;
        RECT 125.000 86.800 130.500 87.100 ;
        RECT 126.500 86.700 126.900 86.800 ;
        RECT 125.700 86.200 126.100 86.300 ;
        RECT 125.700 85.900 128.200 86.200 ;
        RECT 127.800 85.800 128.200 85.900 ;
        RECT 124.600 85.500 127.400 85.600 ;
        RECT 124.600 85.400 127.500 85.500 ;
        RECT 124.600 85.300 129.500 85.400 ;
        RECT 123.800 85.100 124.200 85.200 ;
        RECT 123.000 84.800 124.200 85.100 ;
        RECT 123.000 81.100 123.400 84.800 ;
        RECT 124.600 81.100 125.000 85.300 ;
        RECT 127.100 85.100 129.500 85.300 ;
        RECT 126.200 84.500 128.900 84.800 ;
        RECT 126.200 84.400 126.600 84.500 ;
        RECT 128.500 84.400 128.900 84.500 ;
        RECT 129.200 84.500 129.500 85.100 ;
        RECT 130.200 85.200 130.500 86.800 ;
        RECT 131.000 86.400 131.400 86.500 ;
        RECT 131.000 86.100 132.900 86.400 ;
        RECT 132.500 86.000 132.900 86.100 ;
        RECT 131.700 85.700 132.100 85.800 ;
        RECT 133.400 85.700 133.800 87.400 ;
        RECT 135.800 87.900 136.200 89.900 ;
        RECT 138.200 88.900 138.600 89.900 ;
        RECT 136.500 88.200 136.900 88.600 ;
        RECT 136.600 88.100 137.000 88.200 ;
        RECT 138.200 88.100 138.500 88.900 ;
        RECT 135.000 86.400 135.400 87.200 ;
        RECT 134.200 86.100 134.600 86.200 ;
        RECT 135.800 86.100 136.100 87.900 ;
        RECT 136.600 87.800 138.500 88.100 ;
        RECT 139.000 88.100 139.400 88.600 ;
        RECT 140.600 88.100 141.000 88.200 ;
        RECT 139.000 87.800 141.000 88.100 ;
        RECT 138.200 87.200 138.500 87.800 ;
        RECT 138.200 86.800 138.600 87.200 ;
        RECT 141.400 86.900 141.800 89.900 ;
        RECT 144.600 88.300 145.000 89.900 ;
        RECT 145.400 88.500 145.800 89.900 ;
        RECT 146.200 88.500 146.600 89.900 ;
        RECT 147.000 88.500 147.400 89.900 ;
        RECT 148.600 88.500 149.000 89.900 ;
        RECT 150.200 88.500 150.600 89.900 ;
        RECT 151.000 88.500 151.400 89.900 ;
        RECT 151.800 88.500 152.200 89.900 ;
        RECT 152.600 88.500 153.000 89.900 ;
        RECT 143.700 87.900 145.000 88.300 ;
        RECT 153.400 88.300 153.800 89.900 ;
        RECT 146.700 87.900 149.000 88.200 ;
        RECT 143.700 87.600 144.100 87.900 ;
        RECT 142.600 87.200 144.100 87.600 ;
        RECT 136.600 86.100 137.000 86.200 ;
        RECT 134.200 85.800 135.000 86.100 ;
        RECT 135.800 85.800 137.000 86.100 ;
        RECT 131.700 85.400 133.800 85.700 ;
        RECT 134.600 85.600 135.000 85.800 ;
        RECT 130.200 84.900 131.400 85.200 ;
        RECT 129.900 84.500 130.300 84.600 ;
        RECT 129.200 84.200 130.300 84.500 ;
        RECT 131.100 84.400 131.400 84.900 ;
        RECT 131.100 84.000 131.800 84.400 ;
        RECT 127.900 83.700 128.300 83.800 ;
        RECT 129.300 83.700 129.700 83.800 ;
        RECT 126.200 83.100 126.600 83.500 ;
        RECT 127.900 83.400 129.700 83.700 ;
        RECT 129.000 83.100 129.300 83.400 ;
        RECT 131.000 83.100 131.400 83.500 ;
        RECT 126.200 82.800 127.200 83.100 ;
        RECT 126.800 81.100 127.200 82.800 ;
        RECT 129.000 81.100 129.400 83.100 ;
        RECT 131.100 81.100 131.700 83.100 ;
        RECT 133.400 81.100 133.800 85.400 ;
        RECT 136.600 85.100 136.900 85.800 ;
        RECT 137.400 85.400 137.800 86.200 ;
        RECT 138.200 85.100 138.500 86.800 ;
        RECT 141.400 86.500 145.800 86.900 ;
        RECT 146.700 86.700 147.100 87.900 ;
        RECT 148.600 87.800 149.000 87.900 ;
        RECT 149.400 87.800 150.200 88.200 ;
        RECT 151.700 87.800 152.200 88.200 ;
        RECT 153.400 87.900 154.600 88.300 ;
        RECT 147.800 86.800 148.200 87.600 ;
        RECT 148.600 87.400 149.000 87.500 ;
        RECT 148.600 87.100 150.800 87.400 ;
        RECT 150.400 87.000 150.800 87.100 ;
        RECT 134.200 84.800 136.200 85.100 ;
        RECT 134.200 81.100 134.600 84.800 ;
        RECT 135.800 81.100 136.200 84.800 ;
        RECT 136.600 81.100 137.000 85.100 ;
        RECT 137.700 84.700 138.600 85.100 ;
        RECT 137.700 81.100 138.100 84.700 ;
        RECT 141.400 83.700 141.800 86.500 ;
        RECT 146.100 86.300 147.100 86.700 ;
        RECT 149.000 86.300 150.600 86.700 ;
        RECT 151.800 86.400 152.200 87.800 ;
        RECT 154.200 87.600 154.600 87.900 ;
        RECT 154.200 87.300 155.100 87.600 ;
        RECT 154.700 86.700 155.100 87.300 ;
        RECT 156.600 87.300 157.000 89.900 ;
        RECT 157.400 88.000 157.800 89.900 ;
        RECT 157.400 87.600 157.900 88.000 ;
        RECT 156.600 87.000 157.200 87.300 ;
        RECT 154.700 86.300 156.600 86.700 ;
        RECT 156.900 86.000 157.200 87.000 ;
        RECT 156.800 85.700 157.200 86.000 ;
        RECT 156.800 84.800 157.100 85.700 ;
        RECT 157.500 85.400 157.900 87.600 ;
        RECT 160.600 87.900 161.000 89.900 ;
        RECT 163.000 88.900 163.400 89.900 ;
        RECT 161.300 88.200 161.700 88.600 ;
        RECT 161.400 88.100 161.800 88.200 ;
        RECT 163.000 88.100 163.300 88.900 ;
        RECT 159.800 86.400 160.200 87.200 ;
        RECT 159.000 86.100 159.400 86.200 ;
        RECT 160.600 86.100 160.900 87.900 ;
        RECT 161.400 87.800 163.300 88.100 ;
        RECT 163.000 87.200 163.300 87.800 ;
        RECT 163.800 87.800 164.200 88.600 ;
        RECT 164.600 88.000 165.000 89.900 ;
        RECT 166.200 89.600 168.200 89.900 ;
        RECT 166.200 88.000 166.600 89.600 ;
        RECT 164.600 87.900 166.600 88.000 ;
        RECT 163.800 87.200 164.100 87.800 ;
        RECT 164.700 87.700 166.500 87.900 ;
        RECT 167.000 87.800 167.400 89.300 ;
        RECT 167.800 87.900 168.200 89.600 ;
        RECT 168.600 88.000 169.000 89.900 ;
        RECT 170.200 88.000 170.600 89.900 ;
        RECT 168.600 87.900 170.600 88.000 ;
        RECT 171.000 87.900 171.400 89.900 ;
        RECT 173.400 89.200 173.800 89.900 ;
        RECT 173.400 88.800 173.900 89.200 ;
        RECT 175.000 88.900 175.400 89.900 ;
        RECT 175.000 88.800 175.600 88.900 ;
        RECT 173.600 88.500 175.600 88.800 ;
        RECT 165.000 87.200 165.400 87.400 ;
        RECT 167.100 87.200 167.400 87.800 ;
        RECT 168.700 87.700 170.500 87.900 ;
        RECT 169.000 87.200 169.400 87.400 ;
        RECT 171.000 87.200 171.300 87.900 ;
        RECT 172.600 87.800 173.800 88.200 ;
        RECT 163.000 86.800 163.400 87.200 ;
        RECT 163.800 86.800 164.200 87.200 ;
        RECT 164.600 86.900 165.400 87.200 ;
        RECT 166.200 86.900 167.400 87.200 ;
        RECT 164.600 86.800 165.000 86.900 ;
        RECT 166.200 86.800 166.600 86.900 ;
        RECT 161.400 86.100 161.800 86.200 ;
        RECT 159.000 85.800 159.800 86.100 ;
        RECT 160.600 85.800 161.800 86.100 ;
        RECT 159.400 85.600 159.800 85.800 ;
        RECT 146.200 84.700 146.600 84.800 ;
        RECT 143.900 84.500 146.600 84.700 ;
        RECT 143.500 84.400 146.600 84.500 ;
        RECT 147.100 84.500 151.400 84.800 ;
        RECT 142.200 84.000 143.000 84.400 ;
        RECT 143.500 84.100 144.200 84.400 ;
        RECT 147.100 84.100 147.400 84.500 ;
        RECT 151.000 84.400 151.400 84.500 ;
        RECT 152.600 84.500 157.100 84.800 ;
        RECT 152.600 84.400 153.000 84.500 ;
        RECT 142.700 83.800 143.000 84.000 ;
        RECT 144.500 83.800 147.400 84.100 ;
        RECT 147.700 83.800 149.000 84.200 ;
        RECT 141.400 83.400 142.400 83.700 ;
        RECT 142.700 83.400 144.800 83.800 ;
        RECT 142.100 83.100 142.400 83.400 ;
        RECT 142.100 82.800 142.600 83.100 ;
        RECT 142.200 81.100 142.600 82.800 ;
        RECT 143.800 81.100 144.200 83.400 ;
        RECT 145.400 81.100 145.800 82.500 ;
        RECT 146.200 81.100 146.600 82.500 ;
        RECT 147.000 81.100 147.400 83.500 ;
        RECT 148.600 81.100 149.000 83.500 ;
        RECT 150.200 81.100 150.600 84.200 ;
        RECT 154.200 83.800 155.500 84.200 ;
        RECT 151.800 83.400 153.900 83.800 ;
        RECT 151.000 81.100 151.400 82.500 ;
        RECT 151.800 81.100 152.200 82.500 ;
        RECT 152.600 81.100 153.000 82.500 ;
        RECT 154.200 81.100 154.600 83.800 ;
        RECT 156.800 83.700 157.100 84.500 ;
        RECT 155.800 83.400 157.100 83.700 ;
        RECT 157.400 85.000 157.900 85.400 ;
        RECT 161.400 85.100 161.700 85.800 ;
        RECT 162.200 85.400 162.600 86.200 ;
        RECT 163.000 85.100 163.300 86.800 ;
        RECT 165.400 85.800 165.800 86.600 ;
        RECT 166.200 85.100 166.500 86.800 ;
        RECT 167.000 85.800 167.400 86.600 ;
        RECT 167.800 86.400 168.200 87.200 ;
        RECT 168.600 86.900 169.400 87.200 ;
        RECT 170.100 87.100 171.400 87.200 ;
        RECT 173.400 87.100 174.200 87.200 ;
        RECT 168.600 86.800 169.000 86.900 ;
        RECT 170.100 86.800 174.200 87.100 ;
        RECT 169.400 85.800 169.800 86.600 ;
        RECT 170.100 85.100 170.400 86.800 ;
        RECT 171.000 86.100 171.400 86.200 ;
        RECT 174.200 86.100 175.000 86.200 ;
        RECT 171.000 85.800 175.000 86.100 ;
        RECT 175.300 85.200 175.600 88.500 ;
        RECT 178.200 87.600 178.600 89.900 ;
        RECT 178.200 87.300 179.300 87.600 ;
        RECT 178.200 85.800 178.600 86.600 ;
        RECT 179.000 85.800 179.300 87.300 ;
        RECT 179.000 85.400 179.600 85.800 ;
        RECT 171.000 85.100 171.400 85.200 ;
        RECT 155.800 81.100 156.200 83.400 ;
        RECT 157.400 81.100 157.800 85.000 ;
        RECT 159.000 84.800 161.000 85.100 ;
        RECT 159.000 81.100 159.400 84.800 ;
        RECT 160.600 81.100 161.000 84.800 ;
        RECT 161.400 81.100 161.800 85.100 ;
        RECT 162.500 84.700 163.400 85.100 ;
        RECT 162.500 81.100 162.900 84.700 ;
        RECT 165.900 81.100 166.900 85.100 ;
        RECT 169.900 84.800 170.400 85.100 ;
        RECT 170.700 84.800 171.400 85.100 ;
        RECT 175.300 84.900 177.000 85.200 ;
        RECT 179.000 85.100 179.300 85.400 ;
        RECT 176.600 84.800 177.000 84.900 ;
        RECT 178.200 84.800 179.300 85.100 ;
        RECT 169.900 81.100 170.300 84.800 ;
        RECT 170.700 84.200 171.000 84.800 ;
        RECT 170.600 83.800 171.000 84.200 ;
        RECT 171.900 84.400 173.700 84.700 ;
        RECT 171.900 84.100 172.200 84.400 ;
        RECT 171.800 81.100 172.200 84.100 ;
        RECT 173.400 84.100 173.700 84.400 ;
        RECT 174.300 84.500 176.100 84.600 ;
        RECT 176.600 84.500 176.900 84.800 ;
        RECT 174.300 84.300 176.200 84.500 ;
        RECT 174.300 84.100 174.600 84.300 ;
        RECT 173.400 81.400 173.800 84.100 ;
        RECT 174.200 81.700 174.600 84.100 ;
        RECT 175.000 81.400 175.400 84.000 ;
        RECT 175.800 81.500 176.200 84.300 ;
        RECT 176.600 81.700 177.000 84.500 ;
        RECT 173.400 81.100 175.400 81.400 ;
        RECT 175.900 81.400 176.200 81.500 ;
        RECT 177.400 81.500 177.800 84.500 ;
        RECT 177.400 81.400 177.700 81.500 ;
        RECT 175.900 81.100 177.700 81.400 ;
        RECT 178.200 81.100 178.600 84.800 ;
        RECT 0.600 75.700 1.000 79.900 ;
        RECT 2.800 78.200 3.200 79.900 ;
        RECT 2.200 77.900 3.200 78.200 ;
        RECT 5.000 77.900 5.400 79.900 ;
        RECT 7.100 77.900 7.700 79.900 ;
        RECT 2.200 77.500 2.600 77.900 ;
        RECT 5.000 77.600 5.300 77.900 ;
        RECT 3.900 77.300 5.700 77.600 ;
        RECT 7.000 77.500 7.400 77.900 ;
        RECT 3.900 77.200 4.300 77.300 ;
        RECT 5.300 77.200 5.700 77.300 ;
        RECT 2.200 76.500 2.600 76.600 ;
        RECT 4.500 76.500 4.900 76.600 ;
        RECT 2.200 76.200 4.900 76.500 ;
        RECT 5.200 76.500 6.300 76.800 ;
        RECT 5.200 75.900 5.500 76.500 ;
        RECT 5.900 76.400 6.300 76.500 ;
        RECT 7.100 76.600 7.800 77.000 ;
        RECT 7.100 76.100 7.400 76.600 ;
        RECT 3.100 75.700 5.500 75.900 ;
        RECT 0.600 75.600 5.500 75.700 ;
        RECT 6.200 75.800 7.400 76.100 ;
        RECT 0.600 75.500 3.500 75.600 ;
        RECT 0.600 75.400 3.400 75.500 ;
        RECT 6.200 75.200 6.500 75.800 ;
        RECT 9.400 75.600 9.800 79.900 ;
        RECT 7.700 75.300 9.800 75.600 ;
        RECT 7.700 75.200 8.100 75.300 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 1.700 74.800 4.200 75.100 ;
        RECT 6.200 74.800 6.600 75.200 ;
        RECT 8.500 74.900 8.900 75.000 ;
        RECT 1.700 74.700 2.100 74.800 ;
        RECT 2.500 74.200 2.900 74.300 ;
        RECT 6.200 74.200 6.500 74.800 ;
        RECT 7.000 74.600 8.900 74.900 ;
        RECT 7.000 74.500 7.400 74.600 ;
        RECT 1.000 73.900 6.500 74.200 ;
        RECT 1.000 73.800 1.800 73.900 ;
        RECT 0.600 71.100 1.000 73.500 ;
        RECT 3.100 72.800 3.400 73.900 ;
        RECT 5.900 73.800 6.300 73.900 ;
        RECT 9.400 73.600 9.800 75.300 ;
        RECT 7.900 73.300 9.800 73.600 ;
        RECT 7.900 73.200 8.300 73.300 ;
        RECT 2.200 72.100 2.600 72.500 ;
        RECT 3.000 72.400 3.400 72.800 ;
        RECT 3.900 72.700 4.300 72.800 ;
        RECT 3.900 72.400 5.300 72.700 ;
        RECT 5.000 72.100 5.300 72.400 ;
        RECT 7.000 72.100 7.400 72.500 ;
        RECT 2.200 71.800 3.200 72.100 ;
        RECT 2.800 71.100 3.200 71.800 ;
        RECT 5.000 71.100 5.400 72.100 ;
        RECT 7.000 71.800 7.700 72.100 ;
        RECT 7.100 71.100 7.700 71.800 ;
        RECT 9.400 71.100 9.800 73.300 ;
        RECT 10.200 71.100 10.600 79.900 ;
        RECT 11.800 74.100 12.200 74.200 ;
        RECT 11.000 73.800 12.200 74.100 ;
        RECT 11.000 73.200 11.300 73.800 ;
        RECT 11.800 73.400 12.200 73.800 ;
        RECT 11.000 72.400 11.400 73.200 ;
        RECT 12.600 73.100 13.000 79.900 ;
        RECT 13.400 75.800 13.800 76.600 ;
        RECT 15.000 75.100 15.400 79.900 ;
        RECT 17.700 76.400 18.100 79.900 ;
        RECT 19.800 77.500 20.200 79.500 ;
        RECT 17.300 76.100 18.100 76.400 ;
        RECT 16.600 75.100 17.000 75.600 ;
        RECT 15.000 74.800 17.000 75.100 ;
        RECT 12.600 72.800 13.500 73.100 ;
        RECT 13.100 71.100 13.500 72.800 ;
        RECT 14.200 72.400 14.600 73.200 ;
        RECT 15.000 71.100 15.400 74.800 ;
        RECT 17.300 74.200 17.600 76.100 ;
        RECT 19.900 75.800 20.200 77.500 ;
        RECT 18.300 75.500 20.200 75.800 ;
        RECT 18.300 74.500 18.600 75.500 ;
        RECT 15.800 74.100 16.200 74.200 ;
        RECT 16.600 74.100 17.600 74.200 ;
        RECT 17.900 74.100 18.600 74.500 ;
        RECT 19.000 74.400 19.400 75.200 ;
        RECT 19.800 74.400 20.200 75.200 ;
        RECT 15.800 73.800 17.600 74.100 ;
        RECT 17.300 73.500 17.600 73.800 ;
        RECT 18.100 73.900 18.600 74.100 ;
        RECT 18.100 73.600 20.200 73.900 ;
        RECT 17.300 73.300 17.700 73.500 ;
        RECT 17.300 73.000 18.100 73.300 ;
        RECT 17.700 71.500 18.100 73.000 ;
        RECT 19.900 72.500 20.200 73.600 ;
        RECT 20.600 73.400 21.000 74.200 ;
        RECT 21.400 73.100 21.800 79.900 ;
        RECT 23.800 77.900 24.200 79.900 ;
        RECT 23.900 77.800 24.200 77.900 ;
        RECT 25.400 77.900 25.800 79.900 ;
        RECT 25.400 77.800 25.700 77.900 ;
        RECT 23.900 77.500 25.700 77.800 ;
        RECT 23.000 77.100 23.400 77.200 ;
        RECT 22.200 76.800 23.400 77.100 ;
        RECT 22.200 75.800 22.600 76.800 ;
        RECT 24.600 76.400 25.000 77.200 ;
        RECT 25.400 76.200 25.700 77.500 ;
        RECT 23.000 75.400 23.400 76.200 ;
        RECT 25.400 75.800 25.800 76.200 ;
        RECT 23.800 74.800 24.600 75.200 ;
        RECT 25.400 74.200 25.700 75.800 ;
        RECT 26.200 75.700 26.600 79.900 ;
        RECT 28.400 78.200 28.800 79.900 ;
        RECT 27.800 77.900 28.800 78.200 ;
        RECT 30.600 77.900 31.000 79.900 ;
        RECT 32.700 77.900 33.300 79.900 ;
        RECT 27.800 77.500 28.200 77.900 ;
        RECT 30.600 77.600 30.900 77.900 ;
        RECT 29.500 77.300 31.300 77.600 ;
        RECT 32.600 77.500 33.000 77.900 ;
        RECT 29.500 77.200 29.900 77.300 ;
        RECT 30.900 77.200 31.300 77.300 ;
        RECT 27.800 76.500 28.200 76.600 ;
        RECT 30.100 76.500 30.500 76.600 ;
        RECT 27.800 76.200 30.500 76.500 ;
        RECT 30.800 76.500 31.900 76.800 ;
        RECT 30.800 75.900 31.100 76.500 ;
        RECT 31.500 76.400 31.900 76.500 ;
        RECT 32.700 76.600 33.400 77.000 ;
        RECT 32.700 76.100 33.000 76.600 ;
        RECT 28.700 75.700 31.100 75.900 ;
        RECT 26.200 75.600 31.100 75.700 ;
        RECT 31.800 75.800 33.000 76.100 ;
        RECT 26.200 75.500 29.100 75.600 ;
        RECT 26.200 75.400 29.000 75.500 ;
        RECT 31.800 75.200 32.100 75.800 ;
        RECT 35.000 75.600 35.400 79.900 ;
        RECT 33.300 75.300 35.400 75.600 ;
        RECT 33.300 75.200 33.700 75.300 ;
        RECT 29.400 75.100 29.800 75.200 ;
        RECT 27.300 74.800 29.800 75.100 ;
        RECT 31.800 74.800 32.200 75.200 ;
        RECT 34.100 74.900 34.500 75.000 ;
        RECT 27.300 74.700 27.700 74.800 ;
        RECT 28.100 74.200 28.500 74.300 ;
        RECT 31.800 74.200 32.100 74.800 ;
        RECT 32.600 74.600 34.500 74.900 ;
        RECT 32.600 74.500 33.000 74.600 ;
        RECT 24.900 74.100 25.700 74.200 ;
        RECT 24.800 73.900 25.700 74.100 ;
        RECT 26.600 73.900 32.100 74.200 ;
        RECT 21.400 72.800 22.300 73.100 ;
        RECT 19.800 71.500 20.200 72.500 ;
        RECT 21.900 71.100 22.300 72.800 ;
        RECT 24.800 71.100 25.200 73.900 ;
        RECT 26.600 73.800 27.400 73.900 ;
        RECT 26.200 71.100 26.600 73.500 ;
        RECT 28.700 72.800 29.000 73.900 ;
        RECT 31.500 73.800 31.900 73.900 ;
        RECT 35.000 73.600 35.400 75.300 ;
        RECT 33.500 73.300 35.400 73.600 ;
        RECT 33.500 73.200 33.900 73.300 ;
        RECT 35.000 73.100 35.400 73.300 ;
        RECT 36.600 75.100 37.000 79.900 ;
        RECT 40.900 76.400 41.300 79.900 ;
        RECT 43.000 77.500 43.400 79.500 ;
        RECT 40.500 76.100 41.300 76.400 ;
        RECT 39.800 75.100 40.200 75.600 ;
        RECT 36.600 74.800 40.200 75.100 ;
        RECT 35.800 73.100 36.200 73.200 ;
        RECT 35.000 72.800 36.200 73.100 ;
        RECT 27.800 72.100 28.200 72.500 ;
        RECT 28.600 72.400 29.000 72.800 ;
        RECT 29.500 72.700 29.900 72.800 ;
        RECT 29.500 72.400 30.900 72.700 ;
        RECT 30.600 72.100 30.900 72.400 ;
        RECT 32.600 72.100 33.000 72.500 ;
        RECT 27.800 71.800 28.800 72.100 ;
        RECT 28.400 71.100 28.800 71.800 ;
        RECT 30.600 71.100 31.000 72.100 ;
        RECT 32.600 71.800 33.300 72.100 ;
        RECT 32.700 71.100 33.300 71.800 ;
        RECT 35.000 71.100 35.400 72.800 ;
        RECT 35.800 72.400 36.200 72.800 ;
        RECT 36.600 71.100 37.000 74.800 ;
        RECT 40.500 74.200 40.800 76.100 ;
        RECT 43.100 75.800 43.400 77.500 ;
        RECT 41.500 75.500 43.400 75.800 ;
        RECT 41.500 74.500 41.800 75.500 ;
        RECT 37.400 74.100 37.800 74.200 ;
        RECT 39.800 74.100 40.800 74.200 ;
        RECT 41.100 74.100 41.800 74.500 ;
        RECT 42.200 74.400 42.600 75.200 ;
        RECT 43.000 74.400 43.400 75.200 ;
        RECT 37.400 73.800 40.800 74.100 ;
        RECT 40.500 73.500 40.800 73.800 ;
        RECT 41.300 73.900 41.800 74.100 ;
        RECT 41.300 73.600 43.400 73.900 ;
        RECT 40.500 73.300 40.900 73.500 ;
        RECT 40.500 73.000 41.300 73.300 ;
        RECT 40.900 71.500 41.300 73.000 ;
        RECT 43.100 72.500 43.400 73.600 ;
        RECT 43.800 73.400 44.200 74.200 ;
        RECT 44.600 73.100 45.000 79.900 ;
        RECT 45.400 75.800 45.800 76.600 ;
        RECT 46.200 75.700 46.600 79.900 ;
        RECT 48.400 78.200 48.800 79.900 ;
        RECT 47.800 77.900 48.800 78.200 ;
        RECT 50.600 77.900 51.000 79.900 ;
        RECT 52.700 77.900 53.300 79.900 ;
        RECT 47.800 77.500 48.200 77.900 ;
        RECT 50.600 77.600 50.900 77.900 ;
        RECT 49.500 77.300 51.300 77.600 ;
        RECT 52.600 77.500 53.000 77.900 ;
        RECT 49.500 77.200 49.900 77.300 ;
        RECT 50.900 77.200 51.300 77.300 ;
        RECT 47.800 76.500 48.200 76.600 ;
        RECT 50.100 76.500 50.500 76.600 ;
        RECT 47.800 76.200 50.500 76.500 ;
        RECT 50.800 76.500 51.900 76.800 ;
        RECT 50.800 75.900 51.100 76.500 ;
        RECT 51.500 76.400 51.900 76.500 ;
        RECT 52.700 76.600 53.400 77.000 ;
        RECT 52.700 76.100 53.000 76.600 ;
        RECT 48.700 75.700 51.100 75.900 ;
        RECT 46.200 75.600 51.100 75.700 ;
        RECT 51.800 75.800 53.000 76.100 ;
        RECT 46.200 75.500 49.100 75.600 ;
        RECT 46.200 75.400 49.000 75.500 ;
        RECT 49.400 75.100 49.800 75.200 ;
        RECT 47.300 74.800 49.800 75.100 ;
        RECT 47.300 74.700 47.700 74.800 ;
        RECT 48.100 74.200 48.500 74.300 ;
        RECT 51.800 74.200 52.100 75.800 ;
        RECT 55.000 75.600 55.400 79.900 ;
        RECT 55.800 75.800 56.200 76.600 ;
        RECT 53.300 75.300 55.400 75.600 ;
        RECT 53.300 75.200 53.700 75.300 ;
        RECT 54.100 74.900 54.500 75.000 ;
        RECT 52.600 74.600 54.500 74.900 ;
        RECT 52.600 74.500 53.000 74.600 ;
        RECT 46.600 73.900 52.100 74.200 ;
        RECT 46.600 73.800 47.400 73.900 ;
        RECT 44.600 72.800 45.500 73.100 ;
        RECT 43.000 71.500 43.400 72.500 ;
        RECT 45.100 71.100 45.500 72.800 ;
        RECT 46.200 71.100 46.600 73.500 ;
        RECT 48.700 72.800 49.000 73.900 ;
        RECT 51.500 73.800 51.900 73.900 ;
        RECT 55.000 73.600 55.400 75.300 ;
        RECT 53.500 73.300 55.400 73.600 ;
        RECT 53.500 73.200 53.900 73.300 ;
        RECT 47.800 72.100 48.200 72.500 ;
        RECT 48.600 72.400 49.000 72.800 ;
        RECT 49.500 72.700 49.900 72.800 ;
        RECT 49.500 72.400 50.900 72.700 ;
        RECT 50.600 72.100 50.900 72.400 ;
        RECT 52.600 72.100 53.000 72.500 ;
        RECT 47.800 71.800 48.800 72.100 ;
        RECT 48.400 71.100 48.800 71.800 ;
        RECT 50.600 71.100 51.000 72.100 ;
        RECT 52.600 71.800 53.300 72.100 ;
        RECT 52.700 71.100 53.300 71.800 ;
        RECT 55.000 71.100 55.400 73.300 ;
        RECT 56.600 73.100 57.000 79.900 ;
        RECT 57.400 77.100 57.800 77.200 ;
        RECT 58.200 77.100 58.600 79.900 ;
        RECT 60.300 77.900 60.900 79.900 ;
        RECT 62.600 77.900 63.000 79.900 ;
        RECT 64.800 78.200 65.200 79.900 ;
        RECT 64.800 77.900 65.800 78.200 ;
        RECT 60.600 77.500 61.000 77.900 ;
        RECT 62.700 77.600 63.000 77.900 ;
        RECT 62.300 77.300 64.100 77.600 ;
        RECT 65.400 77.500 65.800 77.900 ;
        RECT 62.300 77.200 62.700 77.300 ;
        RECT 63.700 77.200 64.100 77.300 ;
        RECT 57.400 76.800 58.600 77.100 ;
        RECT 58.200 75.600 58.600 76.800 ;
        RECT 60.200 76.600 60.900 77.000 ;
        RECT 60.600 76.100 60.900 76.600 ;
        RECT 61.700 76.500 62.800 76.800 ;
        RECT 61.700 76.400 62.100 76.500 ;
        RECT 60.600 75.800 61.800 76.100 ;
        RECT 58.200 75.300 60.300 75.600 ;
        RECT 57.400 73.400 57.800 74.200 ;
        RECT 58.200 73.600 58.600 75.300 ;
        RECT 59.900 75.200 60.300 75.300 ;
        RECT 61.500 75.200 61.800 75.800 ;
        RECT 62.500 75.900 62.800 76.500 ;
        RECT 63.100 76.500 63.500 76.600 ;
        RECT 65.400 76.500 65.800 76.600 ;
        RECT 63.100 76.200 65.800 76.500 ;
        RECT 62.500 75.700 64.900 75.900 ;
        RECT 67.000 75.700 67.400 79.900 ;
        RECT 62.500 75.600 67.400 75.700 ;
        RECT 64.500 75.500 67.400 75.600 ;
        RECT 64.600 75.400 67.400 75.500 ;
        RECT 59.100 74.900 59.500 75.000 ;
        RECT 59.100 74.600 61.000 74.900 ;
        RECT 61.400 74.800 61.800 75.200 ;
        RECT 63.000 75.100 63.400 75.200 ;
        RECT 63.800 75.100 64.200 75.200 ;
        RECT 68.600 75.100 69.000 79.900 ;
        RECT 71.300 76.400 71.700 79.900 ;
        RECT 73.400 77.500 73.800 79.500 ;
        RECT 74.200 77.900 74.600 79.900 ;
        RECT 70.900 76.100 71.700 76.400 ;
        RECT 70.200 75.100 70.600 75.600 ;
        RECT 63.000 74.800 66.300 75.100 ;
        RECT 60.600 74.500 61.000 74.600 ;
        RECT 61.500 74.200 61.800 74.800 ;
        RECT 65.900 74.700 66.300 74.800 ;
        RECT 68.600 74.800 70.600 75.100 ;
        RECT 65.100 74.200 65.500 74.300 ;
        RECT 61.500 73.900 67.000 74.200 ;
        RECT 61.700 73.800 62.100 73.900 ;
        RECT 56.100 72.800 57.000 73.100 ;
        RECT 58.200 73.300 60.100 73.600 ;
        RECT 56.100 72.200 56.500 72.800 ;
        RECT 55.800 71.800 56.500 72.200 ;
        RECT 56.100 71.100 56.500 71.800 ;
        RECT 58.200 71.100 58.600 73.300 ;
        RECT 59.700 73.200 60.100 73.300 ;
        RECT 64.600 73.200 64.900 73.900 ;
        RECT 66.200 73.800 67.000 73.900 ;
        RECT 63.700 72.700 64.100 72.800 ;
        RECT 60.600 72.100 61.000 72.500 ;
        RECT 62.700 72.400 64.100 72.700 ;
        RECT 64.600 72.400 65.000 73.200 ;
        RECT 62.700 72.100 63.000 72.400 ;
        RECT 65.400 72.100 65.800 72.500 ;
        RECT 60.300 71.800 61.000 72.100 ;
        RECT 60.300 71.100 60.900 71.800 ;
        RECT 62.600 71.100 63.000 72.100 ;
        RECT 64.800 71.800 65.800 72.100 ;
        RECT 64.800 71.100 65.200 71.800 ;
        RECT 67.000 71.100 67.400 73.500 ;
        RECT 67.800 72.400 68.200 73.200 ;
        RECT 68.600 71.100 69.000 74.800 ;
        RECT 70.900 74.200 71.200 76.100 ;
        RECT 73.500 75.800 73.800 77.500 ;
        RECT 74.300 77.800 74.600 77.900 ;
        RECT 75.800 77.900 76.200 79.900 ;
        RECT 75.800 77.800 76.100 77.900 ;
        RECT 74.300 77.500 76.100 77.800 ;
        RECT 74.300 76.200 74.600 77.500 ;
        RECT 75.000 77.100 75.400 77.200 ;
        RECT 76.600 77.100 77.000 77.200 ;
        RECT 77.400 77.100 77.800 79.900 ;
        RECT 75.000 76.800 77.800 77.100 ;
        RECT 75.000 76.400 75.400 76.800 ;
        RECT 74.200 75.800 74.600 76.200 ;
        RECT 71.900 75.500 73.800 75.800 ;
        RECT 71.900 74.500 72.200 75.500 ;
        RECT 70.200 73.800 71.200 74.200 ;
        RECT 71.500 74.100 72.200 74.500 ;
        RECT 72.600 74.400 73.000 75.200 ;
        RECT 73.400 74.400 73.800 75.200 ;
        RECT 70.900 73.500 71.200 73.800 ;
        RECT 71.700 73.900 72.200 74.100 ;
        RECT 74.300 74.200 74.600 75.800 ;
        RECT 75.400 74.800 76.200 75.200 ;
        RECT 76.600 74.800 77.000 76.200 ;
        RECT 74.300 74.100 75.100 74.200 ;
        RECT 74.300 73.900 75.200 74.100 ;
        RECT 71.700 73.600 73.800 73.900 ;
        RECT 70.900 73.300 71.300 73.500 ;
        RECT 70.900 73.000 71.700 73.300 ;
        RECT 71.300 71.500 71.700 73.000 ;
        RECT 73.500 72.500 73.800 73.600 ;
        RECT 73.400 71.500 73.800 72.500 ;
        RECT 74.800 71.100 75.200 73.900 ;
        RECT 77.400 71.100 77.800 76.800 ;
        RECT 78.200 73.400 78.600 74.200 ;
        RECT 79.000 71.100 79.400 79.900 ;
        RECT 80.600 76.200 81.000 79.900 ;
        RECT 82.200 79.600 84.200 79.900 ;
        RECT 82.200 76.200 82.600 79.600 ;
        RECT 80.600 75.900 82.600 76.200 ;
        RECT 83.000 75.900 83.400 79.300 ;
        RECT 83.800 75.900 84.200 79.600 ;
        RECT 83.000 75.600 83.300 75.900 ;
        RECT 86.200 75.600 86.600 79.900 ;
        RECT 88.300 77.900 88.900 79.900 ;
        RECT 90.600 77.900 91.000 79.900 ;
        RECT 92.800 78.200 93.200 79.900 ;
        RECT 92.800 77.900 93.800 78.200 ;
        RECT 88.600 77.500 89.000 77.900 ;
        RECT 90.700 77.600 91.000 77.900 ;
        RECT 90.300 77.300 92.100 77.600 ;
        RECT 93.400 77.500 93.800 77.900 ;
        RECT 90.300 77.200 90.700 77.300 ;
        RECT 91.700 77.200 92.100 77.300 ;
        RECT 88.200 76.600 88.900 77.000 ;
        RECT 88.600 76.100 88.900 76.600 ;
        RECT 89.700 76.500 90.800 76.800 ;
        RECT 89.700 76.400 90.100 76.500 ;
        RECT 88.600 75.800 89.800 76.100 ;
        RECT 81.000 75.200 81.400 75.400 ;
        RECT 82.300 75.300 83.300 75.600 ;
        RECT 82.300 75.200 82.600 75.300 ;
        RECT 80.600 74.900 81.400 75.200 ;
        RECT 80.600 74.800 81.000 74.900 ;
        RECT 82.200 74.800 82.600 75.200 ;
        RECT 83.800 74.800 84.200 75.600 ;
        RECT 86.200 75.300 88.300 75.600 ;
        RECT 81.400 74.100 81.800 74.600 ;
        RECT 79.800 73.800 81.800 74.100 ;
        RECT 79.800 73.200 80.100 73.800 ;
        RECT 79.800 72.400 80.200 73.200 ;
        RECT 82.300 73.100 82.600 74.800 ;
        RECT 82.900 74.400 83.300 74.800 ;
        RECT 83.000 74.200 83.300 74.400 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 86.200 73.600 86.600 75.300 ;
        RECT 87.900 75.200 88.300 75.300 ;
        RECT 87.100 74.900 87.500 75.000 ;
        RECT 87.100 74.600 89.000 74.900 ;
        RECT 88.600 74.500 89.000 74.600 ;
        RECT 89.500 74.200 89.800 75.800 ;
        RECT 90.500 75.900 90.800 76.500 ;
        RECT 91.100 76.500 91.500 76.600 ;
        RECT 93.400 76.500 93.800 76.600 ;
        RECT 91.100 76.200 93.800 76.500 ;
        RECT 90.500 75.700 92.900 75.900 ;
        RECT 95.000 75.700 95.400 79.900 ;
        RECT 90.500 75.600 95.400 75.700 ;
        RECT 92.500 75.500 95.400 75.600 ;
        RECT 92.600 75.400 95.400 75.500 ;
        RECT 91.000 75.100 91.400 75.200 ;
        RECT 91.800 75.100 92.200 75.200 ;
        RECT 91.000 74.800 94.300 75.100 ;
        RECT 93.900 74.700 94.300 74.800 ;
        RECT 93.100 74.200 93.500 74.300 ;
        RECT 89.500 73.900 95.000 74.200 ;
        RECT 89.700 73.800 90.100 73.900 ;
        RECT 92.600 73.800 93.000 73.900 ;
        RECT 94.200 73.800 95.000 73.900 ;
        RECT 86.200 73.300 88.100 73.600 ;
        RECT 82.100 71.100 82.900 73.100 ;
        RECT 86.200 71.100 86.600 73.300 ;
        RECT 87.700 73.200 88.100 73.300 ;
        RECT 92.600 72.800 92.900 73.800 ;
        RECT 91.700 72.700 92.100 72.800 ;
        RECT 88.600 72.100 89.000 72.500 ;
        RECT 90.700 72.400 92.100 72.700 ;
        RECT 92.600 72.400 93.000 72.800 ;
        RECT 90.700 72.100 91.000 72.400 ;
        RECT 93.400 72.100 93.800 72.500 ;
        RECT 88.300 71.800 89.000 72.100 ;
        RECT 88.300 71.100 88.900 71.800 ;
        RECT 90.600 71.100 91.000 72.100 ;
        RECT 92.800 71.800 93.800 72.100 ;
        RECT 92.800 71.100 93.200 71.800 ;
        RECT 95.000 71.100 95.400 73.500 ;
        RECT 95.800 73.400 96.200 74.200 ;
        RECT 96.600 73.100 97.000 79.900 ;
        RECT 97.400 75.800 97.800 76.600 ;
        RECT 98.200 74.100 98.600 74.200 ;
        RECT 99.000 74.100 99.400 79.900 ;
        RECT 100.900 79.200 101.300 79.900 ;
        RECT 100.600 78.800 101.300 79.200 ;
        RECT 100.900 76.300 101.300 78.800 ;
        RECT 104.300 76.300 104.700 79.900 ;
        RECT 100.900 75.900 101.800 76.300 ;
        RECT 103.800 75.900 104.700 76.300 ;
        RECT 105.400 77.500 105.800 79.500 ;
        RECT 100.600 74.800 101.000 75.600 ;
        RECT 101.400 74.200 101.700 75.900 ;
        RECT 103.900 74.200 104.200 75.900 ;
        RECT 105.400 75.800 105.700 77.500 ;
        RECT 107.500 76.400 107.900 79.900 ;
        RECT 107.500 76.100 108.300 76.400 ;
        RECT 104.600 74.800 105.000 75.600 ;
        RECT 105.400 75.500 107.300 75.800 ;
        RECT 105.400 74.400 105.800 75.200 ;
        RECT 106.200 74.400 106.600 75.200 ;
        RECT 107.000 74.500 107.300 75.500 ;
        RECT 98.200 73.800 99.400 74.100 ;
        RECT 96.600 72.800 97.500 73.100 ;
        RECT 97.100 72.200 97.500 72.800 ;
        RECT 97.100 71.800 97.800 72.200 ;
        RECT 97.100 71.100 97.500 71.800 ;
        RECT 99.000 71.100 99.400 73.800 ;
        RECT 99.800 74.100 100.200 74.200 ;
        RECT 100.600 74.100 101.000 74.200 ;
        RECT 99.800 73.800 101.000 74.100 ;
        RECT 101.400 73.800 101.800 74.200 ;
        RECT 103.800 73.800 104.200 74.200 ;
        RECT 107.000 74.100 107.700 74.500 ;
        RECT 108.000 74.200 108.300 76.100 ;
        RECT 111.500 76.200 111.900 79.900 ;
        RECT 112.200 76.800 112.600 77.200 ;
        RECT 112.300 76.200 112.600 76.800 ;
        RECT 111.500 75.900 112.000 76.200 ;
        RECT 112.300 75.900 113.000 76.200 ;
        RECT 108.600 74.800 109.000 75.600 ;
        RECT 111.000 74.400 111.400 75.200 ;
        RECT 111.700 74.200 112.000 75.900 ;
        RECT 112.600 75.800 113.000 75.900 ;
        RECT 107.000 73.900 107.500 74.100 ;
        RECT 99.800 73.400 100.200 73.800 ;
        RECT 101.400 72.200 101.700 73.800 ;
        RECT 102.200 73.100 102.600 73.200 ;
        RECT 103.000 73.100 103.400 73.200 ;
        RECT 103.900 73.100 104.200 73.800 ;
        RECT 105.400 73.600 107.500 73.900 ;
        RECT 108.000 73.800 109.000 74.200 ;
        RECT 110.200 74.100 110.600 74.200 ;
        RECT 110.200 73.800 111.000 74.100 ;
        RECT 111.700 73.800 113.000 74.200 ;
        RECT 104.600 73.100 105.000 73.200 ;
        RECT 102.200 72.800 103.400 73.100 ;
        RECT 103.800 72.800 105.000 73.100 ;
        RECT 102.200 72.400 102.600 72.800 ;
        RECT 103.000 72.400 103.400 72.800 ;
        RECT 101.400 71.100 101.800 72.200 ;
        RECT 103.900 72.100 104.200 72.800 ;
        RECT 103.800 71.100 104.200 72.100 ;
        RECT 105.400 72.500 105.700 73.600 ;
        RECT 108.000 73.500 108.300 73.800 ;
        RECT 110.600 73.600 111.000 73.800 ;
        RECT 107.900 73.300 108.300 73.500 ;
        RECT 107.500 73.000 108.300 73.300 ;
        RECT 110.300 73.100 112.100 73.300 ;
        RECT 112.600 73.100 112.900 73.800 ;
        RECT 110.200 73.000 112.200 73.100 ;
        RECT 105.400 71.500 105.800 72.500 ;
        RECT 107.500 72.200 107.900 73.000 ;
        RECT 107.500 71.800 108.200 72.200 ;
        RECT 107.500 71.500 107.900 71.800 ;
        RECT 110.200 71.100 110.600 73.000 ;
        RECT 111.800 71.100 112.200 73.000 ;
        RECT 112.600 71.100 113.000 73.100 ;
        RECT 113.400 71.100 113.800 79.900 ;
        RECT 115.100 79.600 116.900 79.900 ;
        RECT 115.100 79.500 115.400 79.600 ;
        RECT 115.000 76.500 115.400 79.500 ;
        RECT 116.600 79.500 116.900 79.600 ;
        RECT 117.400 79.600 119.400 79.900 ;
        RECT 115.800 76.500 116.200 79.300 ;
        RECT 116.600 76.700 117.000 79.500 ;
        RECT 117.400 77.000 117.800 79.600 ;
        RECT 118.200 76.900 118.600 79.300 ;
        RECT 119.000 76.900 119.400 79.600 ;
        RECT 118.200 76.700 118.500 76.900 ;
        RECT 116.600 76.500 118.500 76.700 ;
        RECT 115.900 76.200 116.200 76.500 ;
        RECT 116.700 76.400 118.500 76.500 ;
        RECT 119.100 76.600 119.400 76.900 ;
        RECT 120.600 76.900 121.000 79.900 ;
        RECT 120.600 76.600 120.900 76.900 ;
        RECT 119.100 76.300 120.900 76.600 ;
        RECT 115.800 76.100 116.200 76.200 ;
        RECT 115.800 75.800 117.500 76.100 ;
        RECT 122.700 75.900 123.700 79.900 ;
        RECT 125.400 77.500 125.800 79.500 ;
        RECT 114.200 74.100 114.600 74.200 ;
        RECT 115.800 74.100 116.200 74.200 ;
        RECT 114.200 73.800 116.200 74.100 ;
        RECT 114.200 73.100 114.600 73.200 ;
        RECT 115.800 73.100 116.200 73.200 ;
        RECT 114.200 72.800 116.200 73.100 ;
        RECT 114.200 72.400 114.600 72.800 ;
        RECT 117.200 72.500 117.500 75.800 ;
        RECT 117.800 74.800 118.600 75.200 ;
        RECT 118.200 73.800 119.400 74.200 ;
        RECT 121.400 73.800 121.800 74.600 ;
        RECT 122.200 74.400 122.600 75.200 ;
        RECT 123.100 74.200 123.400 75.900 ;
        RECT 125.400 75.800 125.700 77.500 ;
        RECT 127.500 76.400 127.900 79.900 ;
        RECT 127.500 76.100 128.300 76.400 ;
        RECT 125.400 75.500 127.300 75.800 ;
        RECT 123.800 74.400 124.200 75.200 ;
        RECT 125.400 74.400 125.800 75.200 ;
        RECT 126.200 74.400 126.600 75.200 ;
        RECT 127.000 74.500 127.300 75.500 ;
        RECT 123.000 74.100 123.400 74.200 ;
        RECT 124.600 74.100 125.000 74.200 ;
        RECT 122.200 73.800 123.400 74.100 ;
        RECT 124.200 73.800 125.000 74.100 ;
        RECT 127.000 74.100 127.700 74.500 ;
        RECT 128.000 74.200 128.300 76.100 ;
        RECT 128.600 75.100 129.000 75.600 ;
        RECT 130.200 75.100 130.600 79.900 ;
        RECT 133.700 79.200 134.100 79.900 ;
        RECT 133.400 78.800 134.100 79.200 ;
        RECT 133.700 76.400 134.100 78.800 ;
        RECT 135.800 77.500 136.200 79.500 ;
        RECT 133.300 76.100 134.100 76.400 ;
        RECT 128.600 74.800 130.600 75.100 ;
        RECT 132.600 74.800 133.000 75.600 ;
        RECT 128.000 74.100 129.000 74.200 ;
        RECT 129.400 74.100 129.800 74.200 ;
        RECT 127.000 73.900 127.500 74.100 ;
        RECT 119.000 72.800 120.200 73.200 ;
        RECT 122.200 73.100 122.500 73.800 ;
        RECT 124.200 73.600 124.600 73.800 ;
        RECT 125.400 73.600 127.500 73.900 ;
        RECT 128.000 73.800 129.800 74.100 ;
        RECT 123.100 73.100 124.900 73.300 ;
        RECT 117.200 72.200 119.200 72.500 ;
        RECT 117.200 72.100 117.800 72.200 ;
        RECT 117.400 71.100 117.800 72.100 ;
        RECT 118.900 72.100 119.200 72.200 ;
        RECT 118.900 71.800 119.400 72.100 ;
        RECT 119.000 71.100 119.400 71.800 ;
        RECT 121.400 71.400 121.800 73.100 ;
        RECT 122.200 71.700 122.600 73.100 ;
        RECT 123.000 73.000 125.000 73.100 ;
        RECT 123.000 71.400 123.400 73.000 ;
        RECT 121.400 71.100 123.400 71.400 ;
        RECT 124.600 71.100 125.000 73.000 ;
        RECT 125.400 72.500 125.700 73.600 ;
        RECT 128.000 73.500 128.300 73.800 ;
        RECT 127.900 73.300 128.300 73.500 ;
        RECT 127.500 73.000 128.300 73.300 ;
        RECT 125.400 71.500 125.800 72.500 ;
        RECT 127.500 71.500 127.900 73.000 ;
        RECT 130.200 71.100 130.600 74.800 ;
        RECT 133.300 74.200 133.600 76.100 ;
        RECT 135.900 75.800 136.200 77.500 ;
        RECT 134.300 75.500 136.200 75.800 ;
        RECT 138.200 75.600 138.600 79.900 ;
        RECT 140.300 77.900 140.900 79.900 ;
        RECT 142.600 77.900 143.000 79.900 ;
        RECT 144.800 78.200 145.200 79.900 ;
        RECT 144.800 77.900 145.800 78.200 ;
        RECT 140.600 77.500 141.000 77.900 ;
        RECT 142.700 77.600 143.000 77.900 ;
        RECT 142.300 77.300 144.100 77.600 ;
        RECT 145.400 77.500 145.800 77.900 ;
        RECT 142.300 77.200 142.700 77.300 ;
        RECT 143.700 77.200 144.100 77.300 ;
        RECT 140.200 76.600 140.900 77.000 ;
        RECT 140.600 76.100 140.900 76.600 ;
        RECT 141.700 76.500 142.800 76.800 ;
        RECT 141.700 76.400 142.100 76.500 ;
        RECT 140.600 75.800 141.800 76.100 ;
        RECT 134.300 74.500 134.600 75.500 ;
        RECT 138.200 75.300 140.300 75.600 ;
        RECT 132.600 73.800 133.600 74.200 ;
        RECT 133.900 74.100 134.600 74.500 ;
        RECT 135.000 74.400 135.400 75.200 ;
        RECT 135.800 75.100 136.200 75.200 ;
        RECT 137.400 75.100 137.800 75.200 ;
        RECT 135.800 74.800 137.800 75.100 ;
        RECT 135.800 74.400 136.200 74.800 ;
        RECT 133.300 73.500 133.600 73.800 ;
        RECT 134.100 73.900 134.600 74.100 ;
        RECT 134.100 73.600 136.200 73.900 ;
        RECT 133.300 73.300 133.700 73.500 ;
        RECT 131.000 72.400 131.400 73.200 ;
        RECT 133.300 73.000 134.100 73.300 ;
        RECT 133.700 71.500 134.100 73.000 ;
        RECT 135.900 72.500 136.200 73.600 ;
        RECT 135.800 71.500 136.200 72.500 ;
        RECT 138.200 73.600 138.600 75.300 ;
        RECT 139.900 75.200 140.300 75.300 ;
        RECT 139.100 74.900 139.500 75.000 ;
        RECT 139.100 74.600 141.000 74.900 ;
        RECT 140.600 74.500 141.000 74.600 ;
        RECT 141.500 74.200 141.800 75.800 ;
        RECT 142.500 75.900 142.800 76.500 ;
        RECT 143.100 76.500 143.500 76.600 ;
        RECT 145.400 76.500 145.800 76.600 ;
        RECT 143.100 76.200 145.800 76.500 ;
        RECT 142.500 75.700 144.900 75.900 ;
        RECT 147.000 75.700 147.400 79.900 ;
        RECT 148.600 78.200 149.000 79.900 ;
        RECT 148.500 77.900 149.000 78.200 ;
        RECT 148.500 77.600 148.800 77.900 ;
        RECT 150.200 77.600 150.600 79.900 ;
        RECT 151.800 78.500 152.200 79.900 ;
        RECT 152.600 78.500 153.000 79.900 ;
        RECT 142.500 75.600 147.400 75.700 ;
        RECT 144.500 75.500 147.400 75.600 ;
        RECT 144.600 75.400 147.400 75.500 ;
        RECT 147.800 77.300 148.800 77.600 ;
        RECT 143.800 75.100 144.200 75.200 ;
        RECT 143.800 74.800 146.300 75.100 ;
        RECT 145.900 74.700 146.300 74.800 ;
        RECT 147.800 74.500 148.200 77.300 ;
        RECT 149.100 77.200 151.200 77.600 ;
        RECT 153.400 77.500 153.800 79.900 ;
        RECT 155.000 77.500 155.400 79.900 ;
        RECT 149.100 77.000 149.400 77.200 ;
        RECT 148.600 76.600 149.400 77.000 ;
        RECT 150.900 76.900 153.800 77.200 ;
        RECT 149.900 76.600 150.600 76.900 ;
        RECT 149.900 76.500 153.000 76.600 ;
        RECT 150.300 76.300 153.000 76.500 ;
        RECT 152.600 76.200 153.000 76.300 ;
        RECT 153.500 76.500 153.800 76.900 ;
        RECT 154.100 76.800 155.400 77.200 ;
        RECT 156.600 76.800 157.000 79.900 ;
        RECT 157.400 78.500 157.800 79.900 ;
        RECT 158.200 78.500 158.600 79.900 ;
        RECT 159.000 78.500 159.400 79.900 ;
        RECT 158.200 77.200 160.300 77.600 ;
        RECT 160.600 77.200 161.000 79.900 ;
        RECT 162.200 77.600 162.600 79.900 ;
        RECT 162.200 77.300 163.500 77.600 ;
        RECT 160.600 76.800 161.900 77.200 ;
        RECT 157.400 76.500 157.800 76.600 ;
        RECT 153.500 76.200 157.800 76.500 ;
        RECT 159.000 76.500 159.400 76.600 ;
        RECT 163.200 76.500 163.500 77.300 ;
        RECT 159.000 76.200 163.500 76.500 ;
        RECT 163.200 75.300 163.500 76.200 ;
        RECT 163.800 76.000 164.200 79.900 ;
        RECT 165.400 77.500 165.800 79.500 ;
        RECT 163.800 75.600 164.300 76.000 ;
        RECT 163.200 75.000 163.600 75.300 ;
        RECT 145.100 74.200 145.500 74.300 ;
        RECT 141.500 73.900 147.000 74.200 ;
        RECT 141.700 73.800 142.100 73.900 ;
        RECT 138.200 73.300 140.100 73.600 ;
        RECT 138.200 71.100 138.600 73.300 ;
        RECT 139.700 73.200 140.100 73.300 ;
        RECT 144.600 73.200 144.900 73.900 ;
        RECT 146.200 73.800 147.000 73.900 ;
        RECT 147.800 74.100 152.200 74.500 ;
        RECT 152.500 74.300 153.500 74.700 ;
        RECT 155.400 74.300 157.000 74.700 ;
        RECT 143.700 72.700 144.100 72.800 ;
        RECT 140.600 72.100 141.000 72.500 ;
        RECT 142.700 72.400 144.100 72.700 ;
        RECT 144.600 72.400 145.000 73.200 ;
        RECT 142.700 72.100 143.000 72.400 ;
        RECT 145.400 72.100 145.800 72.500 ;
        RECT 140.300 71.800 141.000 72.100 ;
        RECT 140.300 71.100 140.900 71.800 ;
        RECT 142.600 71.100 143.000 72.100 ;
        RECT 144.800 71.800 145.800 72.100 ;
        RECT 144.800 71.100 145.200 71.800 ;
        RECT 147.000 71.100 147.400 73.500 ;
        RECT 147.800 71.100 148.200 74.100 ;
        RECT 149.000 73.400 150.500 73.800 ;
        RECT 150.100 73.100 150.500 73.400 ;
        RECT 153.100 73.100 153.500 74.300 ;
        RECT 154.200 73.400 154.600 74.200 ;
        RECT 156.800 73.900 157.200 74.000 ;
        RECT 155.000 73.600 157.200 73.900 ;
        RECT 155.000 73.500 155.400 73.600 ;
        RECT 158.200 73.200 158.600 74.600 ;
        RECT 161.100 74.300 163.000 74.700 ;
        RECT 161.100 73.700 161.500 74.300 ;
        RECT 163.300 74.000 163.600 75.000 ;
        RECT 155.000 73.100 155.400 73.200 ;
        RECT 150.100 72.700 151.400 73.100 ;
        RECT 153.100 72.800 155.400 73.100 ;
        RECT 155.800 72.800 156.600 73.200 ;
        RECT 158.100 72.800 158.600 73.200 ;
        RECT 160.600 73.400 161.500 73.700 ;
        RECT 163.000 73.700 163.600 74.000 ;
        RECT 160.600 73.100 161.000 73.400 ;
        RECT 151.000 71.100 151.400 72.700 ;
        RECT 159.800 72.700 161.000 73.100 ;
        RECT 151.800 71.100 152.200 72.500 ;
        RECT 152.600 71.100 153.000 72.500 ;
        RECT 153.400 71.100 153.800 72.500 ;
        RECT 155.000 71.100 155.400 72.500 ;
        RECT 156.600 71.100 157.000 72.500 ;
        RECT 157.400 71.100 157.800 72.500 ;
        RECT 158.200 71.100 158.600 72.500 ;
        RECT 159.000 71.100 159.400 72.500 ;
        RECT 159.800 71.100 160.200 72.700 ;
        RECT 163.000 71.100 163.400 73.700 ;
        RECT 163.900 73.400 164.300 75.600 ;
        RECT 165.400 75.800 165.700 77.500 ;
        RECT 167.500 76.400 167.900 79.900 ;
        RECT 167.500 76.100 168.300 76.400 ;
        RECT 165.400 75.500 167.300 75.800 ;
        RECT 165.400 74.400 165.800 75.200 ;
        RECT 166.200 74.400 166.600 75.200 ;
        RECT 167.000 74.500 167.300 75.500 ;
        RECT 167.000 74.100 167.700 74.500 ;
        RECT 168.000 74.200 168.300 76.100 ;
        RECT 170.200 75.600 170.600 79.900 ;
        RECT 172.300 77.900 172.900 79.900 ;
        RECT 174.600 77.900 175.000 79.900 ;
        RECT 176.800 78.200 177.200 79.900 ;
        RECT 176.800 77.900 177.800 78.200 ;
        RECT 172.600 77.500 173.000 77.900 ;
        RECT 174.700 77.600 175.000 77.900 ;
        RECT 174.300 77.300 176.100 77.600 ;
        RECT 177.400 77.500 177.800 77.900 ;
        RECT 174.300 77.200 174.700 77.300 ;
        RECT 175.700 77.200 176.100 77.300 ;
        RECT 172.200 76.600 172.900 77.000 ;
        RECT 172.600 76.100 172.900 76.600 ;
        RECT 173.700 76.500 174.800 76.800 ;
        RECT 173.700 76.400 174.100 76.500 ;
        RECT 172.600 75.800 173.800 76.100 ;
        RECT 168.600 75.100 169.000 75.600 ;
        RECT 170.200 75.300 172.300 75.600 ;
        RECT 169.400 75.100 169.800 75.200 ;
        RECT 168.600 74.800 169.800 75.100 ;
        RECT 167.000 73.900 167.500 74.100 ;
        RECT 163.800 73.000 164.300 73.400 ;
        RECT 165.400 73.600 167.500 73.900 ;
        RECT 168.000 73.800 169.000 74.200 ;
        RECT 163.800 71.100 164.200 73.000 ;
        RECT 165.400 72.500 165.700 73.600 ;
        RECT 168.000 73.500 168.300 73.800 ;
        RECT 167.900 73.300 168.300 73.500 ;
        RECT 167.500 73.000 168.300 73.300 ;
        RECT 170.200 73.600 170.600 75.300 ;
        RECT 171.900 75.200 172.300 75.300 ;
        RECT 171.100 74.900 171.500 75.000 ;
        RECT 171.100 74.600 173.000 74.900 ;
        RECT 172.600 74.500 173.000 74.600 ;
        RECT 173.500 74.200 173.800 75.800 ;
        RECT 174.500 75.900 174.800 76.500 ;
        RECT 175.100 76.500 175.500 76.600 ;
        RECT 177.400 76.500 177.800 76.600 ;
        RECT 175.100 76.200 177.800 76.500 ;
        RECT 174.500 75.700 176.900 75.900 ;
        RECT 179.000 75.700 179.400 79.900 ;
        RECT 174.500 75.600 179.400 75.700 ;
        RECT 176.500 75.500 179.400 75.600 ;
        RECT 176.600 75.400 179.400 75.500 ;
        RECT 175.800 75.100 176.200 75.200 ;
        RECT 175.800 74.800 178.300 75.100 ;
        RECT 177.900 74.700 178.300 74.800 ;
        RECT 177.100 74.200 177.500 74.300 ;
        RECT 173.500 73.900 179.000 74.200 ;
        RECT 173.700 73.800 174.100 73.900 ;
        RECT 175.800 73.800 176.200 73.900 ;
        RECT 170.200 73.300 172.100 73.600 ;
        RECT 165.400 71.500 165.800 72.500 ;
        RECT 167.500 71.500 167.900 73.000 ;
        RECT 170.200 71.100 170.600 73.300 ;
        RECT 171.700 73.200 172.100 73.300 ;
        RECT 176.600 72.800 176.900 73.900 ;
        RECT 178.200 73.800 179.000 73.900 ;
        RECT 175.700 72.700 176.100 72.800 ;
        RECT 172.600 72.100 173.000 72.500 ;
        RECT 174.700 72.400 176.100 72.700 ;
        RECT 176.600 72.400 177.000 72.800 ;
        RECT 174.700 72.100 175.000 72.400 ;
        RECT 177.400 72.100 177.800 72.500 ;
        RECT 172.300 71.800 173.000 72.100 ;
        RECT 172.300 71.100 172.900 71.800 ;
        RECT 174.600 71.100 175.000 72.100 ;
        RECT 176.800 71.800 177.800 72.100 ;
        RECT 176.800 71.100 177.200 71.800 ;
        RECT 179.000 71.100 179.400 73.500 ;
        RECT 1.400 67.600 1.800 69.900 ;
        RECT 3.000 67.600 3.400 69.900 ;
        RECT 1.400 67.200 3.400 67.600 ;
        RECT 3.000 65.800 3.400 67.200 ;
        RECT 4.600 68.500 5.000 69.500 ;
        RECT 4.600 67.400 4.900 68.500 ;
        RECT 6.700 68.000 7.100 69.500 ;
        RECT 6.700 67.700 7.500 68.000 ;
        RECT 7.100 67.500 7.500 67.700 ;
        RECT 4.600 67.100 6.700 67.400 ;
        RECT 6.200 66.900 6.700 67.100 ;
        RECT 7.200 67.200 7.500 67.500 ;
        RECT 9.400 67.700 9.800 69.900 ;
        RECT 11.500 69.200 12.100 69.900 ;
        RECT 11.500 68.900 12.200 69.200 ;
        RECT 13.800 68.900 14.200 69.900 ;
        RECT 16.000 69.200 16.400 69.900 ;
        RECT 16.000 68.900 17.000 69.200 ;
        RECT 11.800 68.500 12.200 68.900 ;
        RECT 13.900 68.600 14.200 68.900 ;
        RECT 13.900 68.300 15.300 68.600 ;
        RECT 14.900 68.200 15.300 68.300 ;
        RECT 15.800 68.200 16.200 68.600 ;
        RECT 16.600 68.500 17.000 68.900 ;
        RECT 10.900 67.700 11.300 67.800 ;
        RECT 9.400 67.400 11.300 67.700 ;
        RECT 4.600 65.800 5.000 66.600 ;
        RECT 5.400 65.800 5.800 66.600 ;
        RECT 6.200 66.500 6.900 66.900 ;
        RECT 7.200 66.800 8.200 67.200 ;
        RECT 1.400 65.400 3.400 65.800 ;
        RECT 6.200 65.500 6.500 66.500 ;
        RECT 1.400 61.100 1.800 65.400 ;
        RECT 3.000 61.100 3.400 65.400 ;
        RECT 4.600 65.200 6.500 65.500 ;
        RECT 4.600 63.500 4.900 65.200 ;
        RECT 7.200 64.900 7.500 66.800 ;
        RECT 7.800 66.100 8.200 66.200 ;
        RECT 8.600 66.100 9.000 66.200 ;
        RECT 7.800 65.800 9.000 66.100 ;
        RECT 7.800 65.400 8.200 65.800 ;
        RECT 9.400 65.700 9.800 67.400 ;
        RECT 15.800 67.200 16.100 68.200 ;
        RECT 18.200 67.500 18.600 69.900 ;
        RECT 19.000 68.500 19.400 69.500 ;
        RECT 19.000 67.400 19.300 68.500 ;
        RECT 21.100 68.000 21.500 69.500 ;
        RECT 24.100 69.200 24.500 69.900 ;
        RECT 23.800 68.800 24.500 69.200 ;
        RECT 24.100 68.200 24.500 68.800 ;
        RECT 21.100 67.700 21.900 68.000 ;
        RECT 24.100 67.900 25.000 68.200 ;
        RECT 21.500 67.500 21.900 67.700 ;
        RECT 12.900 67.100 13.300 67.200 ;
        RECT 15.800 67.100 16.200 67.200 ;
        RECT 17.400 67.100 18.200 67.200 ;
        RECT 19.000 67.100 21.100 67.400 ;
        RECT 12.700 66.800 18.200 67.100 ;
        RECT 20.600 66.900 21.100 67.100 ;
        RECT 21.600 67.200 21.900 67.500 ;
        RECT 21.600 67.100 22.600 67.200 ;
        RECT 23.800 67.100 24.200 67.200 ;
        RECT 11.800 66.400 12.200 66.500 ;
        RECT 10.300 66.100 12.200 66.400 ;
        RECT 10.300 66.000 10.700 66.100 ;
        RECT 11.100 65.700 11.500 65.800 ;
        RECT 9.400 65.400 11.500 65.700 ;
        RECT 6.700 64.600 7.500 64.900 ;
        RECT 4.600 61.500 5.000 63.500 ;
        RECT 6.700 61.100 7.100 64.600 ;
        RECT 9.400 61.100 9.800 65.400 ;
        RECT 12.700 65.200 13.000 66.800 ;
        RECT 16.300 66.700 16.700 66.800 ;
        RECT 17.100 66.200 17.500 66.300 ;
        RECT 15.000 65.900 17.500 66.200 ;
        RECT 15.000 65.800 15.400 65.900 ;
        RECT 19.000 65.800 19.400 66.600 ;
        RECT 19.800 65.800 20.200 66.600 ;
        RECT 20.600 66.500 21.300 66.900 ;
        RECT 21.600 66.800 24.200 67.100 ;
        RECT 15.800 65.500 18.600 65.600 ;
        RECT 20.600 65.500 20.900 66.500 ;
        RECT 15.700 65.400 18.600 65.500 ;
        RECT 11.800 64.900 13.000 65.200 ;
        RECT 13.700 65.300 18.600 65.400 ;
        RECT 13.700 65.100 16.100 65.300 ;
        RECT 11.800 64.400 12.100 64.900 ;
        RECT 11.400 64.000 12.100 64.400 ;
        RECT 12.900 64.500 13.300 64.600 ;
        RECT 13.700 64.500 14.000 65.100 ;
        RECT 12.900 64.200 14.000 64.500 ;
        RECT 14.300 64.500 17.000 64.800 ;
        RECT 14.300 64.400 14.700 64.500 ;
        RECT 16.600 64.400 17.000 64.500 ;
        RECT 13.500 63.700 13.900 63.800 ;
        RECT 14.900 63.700 15.300 63.800 ;
        RECT 11.800 63.100 12.200 63.500 ;
        RECT 13.500 63.400 15.300 63.700 ;
        RECT 13.900 63.100 14.200 63.400 ;
        RECT 16.600 63.100 17.000 63.500 ;
        RECT 11.500 61.100 12.100 63.100 ;
        RECT 13.800 61.100 14.200 63.100 ;
        RECT 16.000 62.800 17.000 63.100 ;
        RECT 16.000 61.100 16.400 62.800 ;
        RECT 18.200 61.100 18.600 65.300 ;
        RECT 19.000 65.200 20.900 65.500 ;
        RECT 19.000 63.500 19.300 65.200 ;
        RECT 21.600 64.900 21.900 66.800 ;
        RECT 22.200 65.400 22.600 66.200 ;
        RECT 21.100 64.600 21.900 64.900 ;
        RECT 19.000 61.500 19.400 63.500 ;
        RECT 21.100 61.100 21.500 64.600 ;
        RECT 23.800 64.400 24.200 65.200 ;
        RECT 24.600 61.100 25.000 67.900 ;
        RECT 25.400 66.800 25.800 67.600 ;
        RECT 26.200 67.100 26.600 69.900 ;
        RECT 27.000 67.800 27.400 68.600 ;
        RECT 27.800 67.700 28.200 69.900 ;
        RECT 29.900 69.200 30.500 69.900 ;
        RECT 29.900 68.900 30.600 69.200 ;
        RECT 32.200 68.900 32.600 69.900 ;
        RECT 34.400 69.200 34.800 69.900 ;
        RECT 34.400 68.900 35.400 69.200 ;
        RECT 30.200 68.500 30.600 68.900 ;
        RECT 32.300 68.600 32.600 68.900 ;
        RECT 32.300 68.300 33.700 68.600 ;
        RECT 33.300 68.200 33.700 68.300 ;
        RECT 34.200 68.200 34.600 68.600 ;
        RECT 35.000 68.500 35.400 68.900 ;
        RECT 29.300 67.700 29.700 67.800 ;
        RECT 27.800 67.400 29.700 67.700 ;
        RECT 27.000 67.100 27.400 67.200 ;
        RECT 26.200 66.800 27.400 67.100 ;
        RECT 26.200 61.100 26.600 66.800 ;
        RECT 27.800 65.700 28.200 67.400 ;
        RECT 31.300 67.100 31.700 67.200 ;
        RECT 34.200 67.100 34.500 68.200 ;
        RECT 36.600 67.500 37.000 69.900 ;
        RECT 39.000 67.700 39.400 69.900 ;
        RECT 41.100 69.200 41.700 69.900 ;
        RECT 41.100 68.900 41.800 69.200 ;
        RECT 43.400 68.900 43.800 69.900 ;
        RECT 45.600 69.200 46.000 69.900 ;
        RECT 45.600 68.900 46.600 69.200 ;
        RECT 41.400 68.500 41.800 68.900 ;
        RECT 43.500 68.600 43.800 68.900 ;
        RECT 43.500 68.300 44.900 68.600 ;
        RECT 44.500 68.200 44.900 68.300 ;
        RECT 45.400 68.200 45.800 68.600 ;
        RECT 46.200 68.500 46.600 68.900 ;
        RECT 40.500 67.700 40.900 67.800 ;
        RECT 39.000 67.400 40.900 67.700 ;
        RECT 35.800 67.100 36.600 67.200 ;
        RECT 38.200 67.100 38.600 67.200 ;
        RECT 31.100 66.800 38.600 67.100 ;
        RECT 30.200 66.400 30.600 66.500 ;
        RECT 28.700 66.100 30.600 66.400 ;
        RECT 31.100 66.100 31.400 66.800 ;
        RECT 34.700 66.700 35.100 66.800 ;
        RECT 35.500 66.200 35.900 66.300 ;
        RECT 31.800 66.100 32.200 66.200 ;
        RECT 28.700 66.000 29.100 66.100 ;
        RECT 31.000 65.800 32.200 66.100 ;
        RECT 33.400 65.900 35.900 66.200 ;
        RECT 33.400 65.800 33.800 65.900 ;
        RECT 29.500 65.700 29.900 65.800 ;
        RECT 27.800 65.400 29.900 65.700 ;
        RECT 27.800 61.100 28.200 65.400 ;
        RECT 31.100 65.200 31.400 65.800 ;
        RECT 39.000 65.700 39.400 67.400 ;
        RECT 42.500 67.100 42.900 67.200 ;
        RECT 45.400 67.100 45.700 68.200 ;
        RECT 47.800 67.500 48.200 69.900 ;
        RECT 50.200 67.900 50.600 69.900 ;
        RECT 52.600 68.900 53.000 69.900 ;
        RECT 55.800 69.200 56.200 69.900 ;
        RECT 55.800 68.900 56.300 69.200 ;
        RECT 50.900 68.200 51.300 68.600 ;
        RECT 50.200 67.200 50.500 67.900 ;
        RECT 51.000 67.800 51.400 68.200 ;
        RECT 51.800 67.800 52.200 68.600 ;
        RECT 47.000 67.100 47.800 67.200 ;
        RECT 42.300 66.800 47.800 67.100 ;
        RECT 48.600 67.100 49.000 67.200 ;
        RECT 49.400 67.100 49.800 67.200 ;
        RECT 48.600 66.800 49.800 67.100 ;
        RECT 41.400 66.400 41.800 66.500 ;
        RECT 39.900 66.100 41.800 66.400 ;
        RECT 42.300 66.200 42.600 66.800 ;
        RECT 45.900 66.700 46.300 66.800 ;
        RECT 49.400 66.400 49.800 66.800 ;
        RECT 50.200 66.800 50.600 67.200 ;
        RECT 51.000 67.100 51.300 67.800 ;
        RECT 52.700 67.200 53.000 68.900 ;
        RECT 56.000 68.800 56.300 68.900 ;
        RECT 57.400 68.900 57.800 69.900 ;
        RECT 61.400 68.900 61.800 69.900 ;
        RECT 57.400 68.800 58.000 68.900 ;
        RECT 56.000 68.500 58.000 68.800 ;
        RECT 55.000 67.800 55.900 68.200 ;
        RECT 52.600 67.100 53.000 67.200 ;
        RECT 51.000 66.800 53.000 67.100 ;
        RECT 54.200 67.100 54.600 67.200 ;
        RECT 55.800 67.100 56.600 67.200 ;
        RECT 54.200 66.800 56.600 67.100 ;
        RECT 45.400 66.200 45.800 66.300 ;
        RECT 46.700 66.200 47.100 66.300 ;
        RECT 39.900 66.000 40.300 66.100 ;
        RECT 42.200 65.800 42.600 66.200 ;
        RECT 44.600 65.900 47.100 66.200 ;
        RECT 48.600 66.100 49.000 66.200 ;
        RECT 50.200 66.100 50.500 66.800 ;
        RECT 51.000 66.100 51.400 66.200 ;
        RECT 44.600 65.800 45.000 65.900 ;
        RECT 48.600 65.800 49.400 66.100 ;
        RECT 50.200 65.800 51.400 66.100 ;
        RECT 40.700 65.700 41.100 65.800 ;
        RECT 34.200 65.500 37.000 65.600 ;
        RECT 34.100 65.400 37.000 65.500 ;
        RECT 30.200 64.900 31.400 65.200 ;
        RECT 32.100 65.300 37.000 65.400 ;
        RECT 32.100 65.100 34.500 65.300 ;
        RECT 30.200 64.400 30.500 64.900 ;
        RECT 29.800 64.000 30.500 64.400 ;
        RECT 31.300 64.500 31.700 64.600 ;
        RECT 32.100 64.500 32.400 65.100 ;
        RECT 31.300 64.200 32.400 64.500 ;
        RECT 32.700 64.500 35.400 64.800 ;
        RECT 32.700 64.400 33.100 64.500 ;
        RECT 35.000 64.400 35.400 64.500 ;
        RECT 31.900 63.700 32.300 63.800 ;
        RECT 33.300 63.700 33.700 63.800 ;
        RECT 30.200 63.100 30.600 63.500 ;
        RECT 31.900 63.400 33.700 63.700 ;
        RECT 32.300 63.100 32.600 63.400 ;
        RECT 35.000 63.100 35.400 63.500 ;
        RECT 29.900 61.100 30.500 63.100 ;
        RECT 32.200 61.100 32.600 63.100 ;
        RECT 34.400 62.800 35.400 63.100 ;
        RECT 34.400 61.100 34.800 62.800 ;
        RECT 36.600 61.100 37.000 65.300 ;
        RECT 39.000 65.400 41.100 65.700 ;
        RECT 39.000 61.100 39.400 65.400 ;
        RECT 42.300 65.200 42.600 65.800 ;
        RECT 49.000 65.600 49.400 65.800 ;
        RECT 45.400 65.500 48.200 65.600 ;
        RECT 45.300 65.400 48.200 65.500 ;
        RECT 41.400 64.900 42.600 65.200 ;
        RECT 43.300 65.300 48.200 65.400 ;
        RECT 43.300 65.100 45.700 65.300 ;
        RECT 41.400 64.400 41.700 64.900 ;
        RECT 41.000 64.000 41.700 64.400 ;
        RECT 42.500 64.500 42.900 64.600 ;
        RECT 43.300 64.500 43.600 65.100 ;
        RECT 42.500 64.200 43.600 64.500 ;
        RECT 43.900 64.500 46.600 64.800 ;
        RECT 43.900 64.400 44.300 64.500 ;
        RECT 46.200 64.400 46.600 64.500 ;
        RECT 43.100 63.700 43.500 63.800 ;
        RECT 44.500 63.700 44.900 63.800 ;
        RECT 41.400 63.100 41.800 63.500 ;
        RECT 43.100 63.400 44.900 63.700 ;
        RECT 43.500 63.100 43.800 63.400 ;
        RECT 46.200 63.100 46.600 63.500 ;
        RECT 41.100 61.100 41.700 63.100 ;
        RECT 43.400 61.100 43.800 63.100 ;
        RECT 45.600 62.800 46.600 63.100 ;
        RECT 45.600 61.100 46.000 62.800 ;
        RECT 47.800 61.100 48.200 65.300 ;
        RECT 51.000 65.100 51.300 65.800 ;
        RECT 52.700 65.100 53.000 66.800 ;
        RECT 53.400 65.400 53.800 66.200 ;
        RECT 56.600 65.800 57.400 66.200 ;
        RECT 57.700 65.200 58.000 68.500 ;
        RECT 59.800 68.100 60.200 68.200 ;
        RECT 60.600 68.100 61.000 68.600 ;
        RECT 61.500 68.100 61.800 68.900 ;
        RECT 63.100 68.200 63.500 68.600 ;
        RECT 63.000 68.100 63.400 68.200 ;
        RECT 59.800 67.800 61.000 68.100 ;
        RECT 61.400 67.800 63.400 68.100 ;
        RECT 63.800 67.900 64.200 69.900 ;
        RECT 61.500 67.200 61.800 67.800 ;
        RECT 61.400 66.800 61.800 67.200 ;
        RECT 59.800 65.800 60.200 66.200 ;
        RECT 57.700 65.100 59.400 65.200 ;
        RECT 59.800 65.100 60.100 65.800 ;
        RECT 61.500 65.100 61.800 66.800 ;
        RECT 62.200 65.400 62.600 66.200 ;
        RECT 63.000 66.100 63.400 66.200 ;
        RECT 63.900 66.100 64.200 67.900 ;
        RECT 64.600 66.400 65.000 67.200 ;
        RECT 65.400 66.100 65.800 66.200 ;
        RECT 66.200 66.100 66.600 66.200 ;
        RECT 63.000 65.800 64.200 66.100 ;
        RECT 65.000 65.800 66.600 66.100 ;
        RECT 63.100 65.100 63.400 65.800 ;
        RECT 65.000 65.600 65.400 65.800 ;
        RECT 48.600 64.800 50.600 65.100 ;
        RECT 48.600 61.100 49.000 64.800 ;
        RECT 50.200 61.100 50.600 64.800 ;
        RECT 51.000 61.100 51.400 65.100 ;
        RECT 52.600 64.700 53.500 65.100 ;
        RECT 57.700 64.900 60.100 65.100 ;
        RECT 59.000 64.800 60.100 64.900 ;
        RECT 53.100 61.100 53.500 64.700 ;
        RECT 54.300 64.400 56.100 64.700 ;
        RECT 54.300 64.100 54.600 64.400 ;
        RECT 54.200 61.100 54.600 64.100 ;
        RECT 55.800 64.100 56.100 64.400 ;
        RECT 56.700 64.500 58.500 64.600 ;
        RECT 59.000 64.500 59.300 64.800 ;
        RECT 61.400 64.700 62.300 65.100 ;
        RECT 56.700 64.300 58.600 64.500 ;
        RECT 56.700 64.100 57.000 64.300 ;
        RECT 55.800 61.400 56.200 64.100 ;
        RECT 56.600 61.700 57.000 64.100 ;
        RECT 57.400 61.400 57.800 64.000 ;
        RECT 58.200 61.500 58.600 64.300 ;
        RECT 59.000 61.700 59.400 64.500 ;
        RECT 55.800 61.100 57.800 61.400 ;
        RECT 58.300 61.400 58.600 61.500 ;
        RECT 59.800 61.500 60.200 64.500 ;
        RECT 59.800 61.400 60.100 61.500 ;
        RECT 58.300 61.100 60.100 61.400 ;
        RECT 61.900 61.100 62.300 64.700 ;
        RECT 63.000 61.100 63.400 65.100 ;
        RECT 63.800 64.800 65.800 65.100 ;
        RECT 63.800 61.100 64.200 64.800 ;
        RECT 65.400 61.100 65.800 64.800 ;
        RECT 67.000 61.100 67.400 69.900 ;
        RECT 67.800 66.800 68.200 67.600 ;
        RECT 68.600 66.800 69.000 67.600 ;
        RECT 69.400 61.100 69.800 69.900 ;
        RECT 70.200 67.500 70.600 69.900 ;
        RECT 72.400 69.200 72.800 69.900 ;
        RECT 71.800 68.900 72.800 69.200 ;
        RECT 74.600 68.900 75.000 69.900 ;
        RECT 76.700 69.200 77.300 69.900 ;
        RECT 76.600 68.900 77.300 69.200 ;
        RECT 71.800 68.500 72.200 68.900 ;
        RECT 74.600 68.600 74.900 68.900 ;
        RECT 72.600 67.800 73.000 68.600 ;
        RECT 73.500 68.300 74.900 68.600 ;
        RECT 76.600 68.500 77.000 68.900 ;
        RECT 73.500 68.200 73.900 68.300 ;
        RECT 79.000 68.100 79.400 69.900 ;
        RECT 79.800 68.100 80.200 68.600 ;
        RECT 79.000 67.800 80.200 68.100 ;
        RECT 70.600 67.100 71.400 67.200 ;
        RECT 72.700 67.100 73.000 67.800 ;
        RECT 77.500 67.700 77.900 67.800 ;
        RECT 79.000 67.700 79.400 67.800 ;
        RECT 77.500 67.400 79.400 67.700 ;
        RECT 75.500 67.100 75.900 67.200 ;
        RECT 70.600 66.800 76.100 67.100 ;
        RECT 72.100 66.700 72.500 66.800 ;
        RECT 71.300 66.200 71.700 66.300 ;
        RECT 71.300 65.900 73.800 66.200 ;
        RECT 73.400 65.800 73.800 65.900 ;
        RECT 70.200 65.500 73.000 65.600 ;
        RECT 70.200 65.400 73.100 65.500 ;
        RECT 70.200 65.300 75.100 65.400 ;
        RECT 70.200 61.100 70.600 65.300 ;
        RECT 72.700 65.100 75.100 65.300 ;
        RECT 71.800 64.500 74.500 64.800 ;
        RECT 71.800 64.400 72.200 64.500 ;
        RECT 74.100 64.400 74.500 64.500 ;
        RECT 74.800 64.500 75.100 65.100 ;
        RECT 75.800 65.200 76.100 66.800 ;
        RECT 76.600 66.400 77.000 66.500 ;
        RECT 76.600 66.100 78.500 66.400 ;
        RECT 78.100 66.000 78.500 66.100 ;
        RECT 77.300 65.700 77.700 65.800 ;
        RECT 79.000 65.700 79.400 67.400 ;
        RECT 77.300 65.400 79.400 65.700 ;
        RECT 75.800 64.900 77.000 65.200 ;
        RECT 75.500 64.500 75.900 64.600 ;
        RECT 74.800 64.200 75.900 64.500 ;
        RECT 76.700 64.400 77.000 64.900 ;
        RECT 76.700 64.000 77.400 64.400 ;
        RECT 73.500 63.700 73.900 63.800 ;
        RECT 74.900 63.700 75.300 63.800 ;
        RECT 71.800 63.100 72.200 63.500 ;
        RECT 73.500 63.400 75.300 63.700 ;
        RECT 74.600 63.100 74.900 63.400 ;
        RECT 76.600 63.100 77.000 63.500 ;
        RECT 71.800 62.800 72.800 63.100 ;
        RECT 72.400 61.100 72.800 62.800 ;
        RECT 74.600 61.100 75.000 63.100 ;
        RECT 76.700 61.100 77.300 63.100 ;
        RECT 79.000 61.100 79.400 65.400 ;
        RECT 80.600 66.100 81.000 69.900 ;
        RECT 83.300 68.000 83.700 69.500 ;
        RECT 85.400 68.500 85.800 69.500 ;
        RECT 87.500 69.200 88.300 69.900 ;
        RECT 87.000 68.800 88.300 69.200 ;
        RECT 91.000 69.100 91.400 69.200 ;
        RECT 91.800 69.100 92.200 69.900 ;
        RECT 91.000 68.800 92.200 69.100 ;
        RECT 93.900 69.200 94.500 69.900 ;
        RECT 93.900 68.900 94.600 69.200 ;
        RECT 96.200 68.900 96.600 69.900 ;
        RECT 98.400 69.200 98.800 69.900 ;
        RECT 98.400 68.900 99.400 69.200 ;
        RECT 82.900 67.700 83.700 68.000 ;
        RECT 82.900 67.500 83.300 67.700 ;
        RECT 82.900 67.200 83.200 67.500 ;
        RECT 85.500 67.400 85.800 68.500 ;
        RECT 87.500 67.900 88.300 68.800 ;
        RECT 81.400 67.100 81.800 67.200 ;
        RECT 82.200 67.100 83.200 67.200 ;
        RECT 81.400 66.800 83.200 67.100 ;
        RECT 83.700 67.100 85.800 67.400 ;
        RECT 86.200 67.100 86.600 67.200 ;
        RECT 87.000 67.100 87.400 67.200 ;
        RECT 83.700 66.900 84.200 67.100 ;
        RECT 82.200 66.100 82.600 66.200 ;
        RECT 80.600 65.800 82.600 66.100 ;
        RECT 80.600 61.100 81.000 65.800 ;
        RECT 82.200 65.400 82.600 65.800 ;
        RECT 82.900 64.900 83.200 66.800 ;
        RECT 83.500 66.500 84.200 66.900 ;
        RECT 86.200 66.800 87.400 67.100 ;
        RECT 87.100 66.600 87.400 66.800 ;
        RECT 83.900 65.500 84.200 66.500 ;
        RECT 84.600 65.800 85.000 66.600 ;
        RECT 85.400 65.800 85.800 66.600 ;
        RECT 87.100 66.200 87.500 66.600 ;
        RECT 87.800 66.200 88.100 67.900 ;
        RECT 91.800 67.700 92.200 68.800 ;
        RECT 94.200 68.500 94.600 68.900 ;
        RECT 96.300 68.600 96.600 68.900 ;
        RECT 96.300 68.300 97.700 68.600 ;
        RECT 97.300 68.200 97.700 68.300 ;
        RECT 98.200 67.800 98.600 68.600 ;
        RECT 99.000 68.500 99.400 68.900 ;
        RECT 93.300 67.700 93.700 67.800 ;
        RECT 91.800 67.400 93.700 67.700 ;
        RECT 88.600 67.100 89.000 67.200 ;
        RECT 91.000 67.100 91.400 67.200 ;
        RECT 88.600 66.800 91.400 67.100 ;
        RECT 88.600 66.400 89.000 66.800 ;
        RECT 83.900 65.200 85.800 65.500 ;
        RECT 86.200 65.400 86.600 66.200 ;
        RECT 87.800 65.800 88.200 66.200 ;
        RECT 89.400 66.100 89.800 66.200 ;
        RECT 89.000 65.800 89.800 66.100 ;
        RECT 87.800 65.700 88.100 65.800 ;
        RECT 87.100 65.400 88.100 65.700 ;
        RECT 89.000 65.600 89.400 65.800 ;
        RECT 91.800 65.700 92.200 67.400 ;
        RECT 95.300 67.100 95.700 67.200 ;
        RECT 98.200 67.100 98.500 67.800 ;
        RECT 100.600 67.500 101.000 69.900 ;
        RECT 101.400 67.800 101.800 68.600 ;
        RECT 99.800 67.100 100.600 67.200 ;
        RECT 95.100 66.800 100.600 67.100 ;
        RECT 94.200 66.400 94.600 66.500 ;
        RECT 92.700 66.100 94.600 66.400 ;
        RECT 92.700 66.000 93.100 66.100 ;
        RECT 93.500 65.700 93.900 65.800 ;
        RECT 91.800 65.400 93.900 65.700 ;
        RECT 82.900 64.600 83.700 64.900 ;
        RECT 83.300 61.100 83.700 64.600 ;
        RECT 85.500 63.500 85.800 65.200 ;
        RECT 87.100 65.100 87.400 65.400 ;
        RECT 85.400 61.500 85.800 63.500 ;
        RECT 86.200 61.400 86.600 65.100 ;
        RECT 87.000 61.700 87.400 65.100 ;
        RECT 87.800 64.800 89.800 65.100 ;
        RECT 87.800 61.400 88.200 64.800 ;
        RECT 86.200 61.100 88.200 61.400 ;
        RECT 89.400 61.100 89.800 64.800 ;
        RECT 91.800 61.100 92.200 65.400 ;
        RECT 95.100 65.200 95.400 66.800 ;
        RECT 98.700 66.700 99.100 66.800 ;
        RECT 98.200 66.200 98.600 66.300 ;
        RECT 99.500 66.200 99.900 66.300 ;
        RECT 97.400 65.900 99.900 66.200 ;
        RECT 102.200 66.100 102.600 69.900 ;
        RECT 104.900 68.000 105.300 69.500 ;
        RECT 107.000 68.500 107.400 69.500 ;
        RECT 104.500 67.700 105.300 68.000 ;
        RECT 104.500 67.500 104.900 67.700 ;
        RECT 104.500 67.200 104.800 67.500 ;
        RECT 107.100 67.400 107.400 68.500 ;
        RECT 107.800 67.500 108.200 69.900 ;
        RECT 110.000 69.200 110.400 69.900 ;
        RECT 109.400 68.900 110.400 69.200 ;
        RECT 112.200 68.900 112.600 69.900 ;
        RECT 114.300 69.200 114.900 69.900 ;
        RECT 114.200 68.900 114.900 69.200 ;
        RECT 109.400 68.500 109.800 68.900 ;
        RECT 112.200 68.600 112.500 68.900 ;
        RECT 110.200 67.800 110.600 68.600 ;
        RECT 111.100 68.300 112.500 68.600 ;
        RECT 114.200 68.500 114.600 68.900 ;
        RECT 111.100 68.200 111.500 68.300 ;
        RECT 103.000 67.100 103.400 67.200 ;
        RECT 103.800 67.100 104.800 67.200 ;
        RECT 103.000 66.800 104.800 67.100 ;
        RECT 105.300 67.100 107.400 67.400 ;
        RECT 108.200 67.100 109.000 67.200 ;
        RECT 110.300 67.100 110.600 67.800 ;
        RECT 115.100 67.700 115.500 67.800 ;
        RECT 116.600 67.700 117.000 69.900 ;
        RECT 118.200 68.800 118.600 69.900 ;
        RECT 117.400 67.800 117.800 68.600 ;
        RECT 115.100 67.400 117.000 67.700 ;
        RECT 113.100 67.100 113.500 67.200 ;
        RECT 105.300 66.900 105.800 67.100 ;
        RECT 103.800 66.100 104.200 66.200 ;
        RECT 97.400 65.800 97.800 65.900 ;
        RECT 102.200 65.800 104.200 66.100 ;
        RECT 98.200 65.500 101.000 65.600 ;
        RECT 98.100 65.400 101.000 65.500 ;
        RECT 94.200 64.900 95.400 65.200 ;
        RECT 96.100 65.300 101.000 65.400 ;
        RECT 96.100 65.100 98.500 65.300 ;
        RECT 94.200 64.400 94.500 64.900 ;
        RECT 93.800 64.000 94.500 64.400 ;
        RECT 95.300 64.500 95.700 64.600 ;
        RECT 96.100 64.500 96.400 65.100 ;
        RECT 95.300 64.200 96.400 64.500 ;
        RECT 96.700 64.500 99.400 64.800 ;
        RECT 96.700 64.400 97.100 64.500 ;
        RECT 99.000 64.400 99.400 64.500 ;
        RECT 95.900 63.700 96.300 63.800 ;
        RECT 97.300 63.700 97.700 63.800 ;
        RECT 94.200 63.100 94.600 63.500 ;
        RECT 95.900 63.400 97.700 63.700 ;
        RECT 96.300 63.100 96.600 63.400 ;
        RECT 99.000 63.100 99.400 63.500 ;
        RECT 93.900 61.100 94.500 63.100 ;
        RECT 96.200 61.100 96.600 63.100 ;
        RECT 98.400 62.800 99.400 63.100 ;
        RECT 98.400 61.100 98.800 62.800 ;
        RECT 100.600 61.100 101.000 65.300 ;
        RECT 102.200 61.100 102.600 65.800 ;
        RECT 103.800 65.400 104.200 65.800 ;
        RECT 104.500 64.900 104.800 66.800 ;
        RECT 105.100 66.500 105.800 66.900 ;
        RECT 108.200 66.800 113.700 67.100 ;
        RECT 109.700 66.700 110.100 66.800 ;
        RECT 105.500 65.500 105.800 66.500 ;
        RECT 106.200 65.800 106.600 66.600 ;
        RECT 107.000 65.800 107.400 66.600 ;
        RECT 108.900 66.200 109.300 66.300 ;
        RECT 108.900 65.900 111.400 66.200 ;
        RECT 111.000 65.800 111.400 65.900 ;
        RECT 107.800 65.500 110.600 65.600 ;
        RECT 105.500 65.200 107.400 65.500 ;
        RECT 104.500 64.600 105.300 64.900 ;
        RECT 104.900 61.100 105.300 64.600 ;
        RECT 107.100 63.500 107.400 65.200 ;
        RECT 107.000 61.500 107.400 63.500 ;
        RECT 107.800 65.400 110.700 65.500 ;
        RECT 107.800 65.300 112.700 65.400 ;
        RECT 107.800 61.100 108.200 65.300 ;
        RECT 110.300 65.100 112.700 65.300 ;
        RECT 109.400 64.500 112.100 64.800 ;
        RECT 109.400 64.400 109.800 64.500 ;
        RECT 111.700 64.400 112.100 64.500 ;
        RECT 112.400 64.500 112.700 65.100 ;
        RECT 113.400 65.200 113.700 66.800 ;
        RECT 114.200 66.400 114.600 66.500 ;
        RECT 114.200 66.100 116.100 66.400 ;
        RECT 115.700 66.000 116.100 66.100 ;
        RECT 114.900 65.700 115.300 65.800 ;
        RECT 116.600 65.700 117.000 67.400 ;
        RECT 118.300 67.200 118.600 68.800 ;
        RECT 118.200 66.800 118.600 67.200 ;
        RECT 119.800 68.500 120.200 69.500 ;
        RECT 119.800 67.400 120.100 68.500 ;
        RECT 121.900 68.000 122.300 69.500 ;
        RECT 121.900 67.700 122.700 68.000 ;
        RECT 122.300 67.500 122.700 67.700 ;
        RECT 124.600 67.500 125.000 69.900 ;
        RECT 126.800 69.200 127.200 69.900 ;
        RECT 126.200 68.900 127.200 69.200 ;
        RECT 129.000 68.900 129.400 69.900 ;
        RECT 131.100 69.200 131.700 69.900 ;
        RECT 131.000 68.900 131.700 69.200 ;
        RECT 126.200 68.500 126.600 68.900 ;
        RECT 129.000 68.600 129.300 68.900 ;
        RECT 127.000 67.800 127.400 68.600 ;
        RECT 127.900 68.300 129.300 68.600 ;
        RECT 131.000 68.500 131.400 68.900 ;
        RECT 127.900 68.200 128.300 68.300 ;
        RECT 133.400 68.100 133.800 69.900 ;
        RECT 134.200 68.100 134.600 68.600 ;
        RECT 133.400 67.800 134.600 68.100 ;
        RECT 119.800 67.100 121.900 67.400 ;
        RECT 114.900 65.400 117.000 65.700 ;
        RECT 113.400 64.900 114.600 65.200 ;
        RECT 113.100 64.500 113.500 64.600 ;
        RECT 112.400 64.200 113.500 64.500 ;
        RECT 114.300 64.400 114.600 64.900 ;
        RECT 114.300 64.000 115.000 64.400 ;
        RECT 111.100 63.700 111.500 63.800 ;
        RECT 112.500 63.700 112.900 63.800 ;
        RECT 109.400 63.100 109.800 63.500 ;
        RECT 111.100 63.400 112.900 63.700 ;
        RECT 112.200 63.100 112.500 63.400 ;
        RECT 114.200 63.100 114.600 63.500 ;
        RECT 109.400 62.800 110.400 63.100 ;
        RECT 110.000 61.100 110.400 62.800 ;
        RECT 112.200 61.100 112.600 63.100 ;
        RECT 114.300 61.100 114.900 63.100 ;
        RECT 116.600 61.100 117.000 65.400 ;
        RECT 118.300 65.100 118.600 66.800 ;
        RECT 121.400 66.900 121.900 67.100 ;
        RECT 122.400 67.200 122.700 67.500 ;
        RECT 119.000 65.400 119.400 66.200 ;
        RECT 119.800 65.800 120.200 66.600 ;
        RECT 120.600 65.800 121.000 66.600 ;
        RECT 121.400 66.500 122.100 66.900 ;
        RECT 122.400 66.800 123.400 67.200 ;
        RECT 125.000 67.100 125.800 67.200 ;
        RECT 127.100 67.100 127.400 67.800 ;
        RECT 131.900 67.700 132.300 67.800 ;
        RECT 133.400 67.700 133.800 67.800 ;
        RECT 131.900 67.400 133.800 67.700 ;
        RECT 129.900 67.100 130.300 67.200 ;
        RECT 125.000 66.800 130.500 67.100 ;
        RECT 121.400 65.500 121.700 66.500 ;
        RECT 119.800 65.200 121.700 65.500 ;
        RECT 118.200 64.700 119.100 65.100 ;
        RECT 118.700 61.100 119.100 64.700 ;
        RECT 119.800 63.500 120.100 65.200 ;
        RECT 122.400 64.900 122.700 66.800 ;
        RECT 126.500 66.700 126.900 66.800 ;
        RECT 125.700 66.200 126.100 66.300 ;
        RECT 127.000 66.200 127.400 66.300 ;
        RECT 123.000 66.100 123.400 66.200 ;
        RECT 123.800 66.100 124.200 66.200 ;
        RECT 123.000 65.800 124.200 66.100 ;
        RECT 125.700 65.900 128.200 66.200 ;
        RECT 127.800 65.800 128.200 65.900 ;
        RECT 123.000 65.400 123.400 65.800 ;
        RECT 124.600 65.500 127.400 65.600 ;
        RECT 124.600 65.400 127.500 65.500 ;
        RECT 121.900 64.600 122.700 64.900 ;
        RECT 124.600 65.300 129.500 65.400 ;
        RECT 119.800 61.500 120.200 63.500 ;
        RECT 121.900 61.100 122.300 64.600 ;
        RECT 124.600 61.100 125.000 65.300 ;
        RECT 127.100 65.100 129.500 65.300 ;
        RECT 126.200 64.500 128.900 64.800 ;
        RECT 126.200 64.400 126.600 64.500 ;
        RECT 128.500 64.400 128.900 64.500 ;
        RECT 129.200 64.500 129.500 65.100 ;
        RECT 130.200 65.200 130.500 66.800 ;
        RECT 131.000 66.400 131.400 66.500 ;
        RECT 131.000 66.100 132.900 66.400 ;
        RECT 132.500 66.000 132.900 66.100 ;
        RECT 131.700 65.700 132.100 65.800 ;
        RECT 133.400 65.700 133.800 67.400 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 135.000 66.100 135.400 69.900 ;
        RECT 135.800 69.600 137.800 69.900 ;
        RECT 135.800 67.900 136.200 69.600 ;
        RECT 136.600 67.900 137.000 69.300 ;
        RECT 137.400 68.000 137.800 69.600 ;
        RECT 139.000 68.000 139.400 69.900 ;
        RECT 137.400 67.900 139.400 68.000 ;
        RECT 141.400 69.600 143.400 69.900 ;
        RECT 141.400 67.900 141.800 69.600 ;
        RECT 142.200 67.900 142.600 69.300 ;
        RECT 143.000 68.000 143.400 69.600 ;
        RECT 144.600 68.000 145.000 69.900 ;
        RECT 147.000 69.200 147.400 69.900 ;
        RECT 147.000 68.800 147.500 69.200 ;
        RECT 148.600 68.900 149.000 69.900 ;
        RECT 148.600 68.800 149.200 68.900 ;
        RECT 147.200 68.500 149.200 68.800 ;
        RECT 143.000 67.900 145.000 68.000 ;
        RECT 136.600 67.200 136.900 67.900 ;
        RECT 137.500 67.700 139.300 67.900 ;
        RECT 138.600 67.200 139.000 67.400 ;
        RECT 142.200 67.200 142.500 67.900 ;
        RECT 143.100 67.700 144.900 67.900 ;
        RECT 146.200 67.800 147.100 68.200 ;
        RECT 144.200 67.200 144.600 67.400 ;
        RECT 135.800 66.400 136.200 67.200 ;
        RECT 136.600 66.900 137.800 67.200 ;
        RECT 138.600 66.900 139.400 67.200 ;
        RECT 137.400 66.800 137.800 66.900 ;
        RECT 139.000 66.800 139.400 66.900 ;
        RECT 134.200 65.800 135.400 66.100 ;
        RECT 136.600 65.800 137.000 66.600 ;
        RECT 131.700 65.400 133.800 65.700 ;
        RECT 130.200 64.900 131.400 65.200 ;
        RECT 129.900 64.500 130.300 64.600 ;
        RECT 129.200 64.200 130.300 64.500 ;
        RECT 131.100 64.400 131.400 64.900 ;
        RECT 131.100 64.000 131.800 64.400 ;
        RECT 127.900 63.700 128.300 63.800 ;
        RECT 129.300 63.700 129.700 63.800 ;
        RECT 126.200 63.100 126.600 63.500 ;
        RECT 127.900 63.400 129.700 63.700 ;
        RECT 129.000 63.100 129.300 63.400 ;
        RECT 131.000 63.100 131.400 63.500 ;
        RECT 126.200 62.800 127.200 63.100 ;
        RECT 126.800 61.100 127.200 62.800 ;
        RECT 129.000 61.100 129.400 63.100 ;
        RECT 131.100 61.100 131.700 63.100 ;
        RECT 133.400 61.100 133.800 65.400 ;
        RECT 135.000 61.100 135.400 65.800 ;
        RECT 137.500 65.100 137.800 66.800 ;
        RECT 138.200 65.800 138.600 66.600 ;
        RECT 141.400 66.400 141.800 67.200 ;
        RECT 142.200 66.900 143.400 67.200 ;
        RECT 144.200 66.900 145.000 67.200 ;
        RECT 143.000 66.800 143.400 66.900 ;
        RECT 144.600 66.800 145.000 66.900 ;
        RECT 147.000 66.800 148.200 67.200 ;
        RECT 142.200 65.800 142.600 66.600 ;
        RECT 143.100 65.200 143.400 66.800 ;
        RECT 143.800 65.800 144.200 66.600 ;
        RECT 147.800 65.800 148.600 66.200 ;
        RECT 148.900 65.200 149.200 68.500 ;
        RECT 153.400 67.900 153.800 69.900 ;
        RECT 154.100 68.200 154.500 68.600 ;
        RECT 150.200 67.100 150.600 67.200 ;
        RECT 151.800 67.100 152.200 67.200 ;
        RECT 150.200 66.800 152.200 67.100 ;
        RECT 152.600 66.400 153.000 67.200 ;
        RECT 151.800 66.100 152.200 66.200 ;
        RECT 153.400 66.100 153.700 67.900 ;
        RECT 154.200 67.800 154.600 68.200 ;
        RECT 155.000 67.900 155.400 69.900 ;
        RECT 155.800 68.000 156.200 69.900 ;
        RECT 157.400 68.000 157.800 69.900 ;
        RECT 163.000 69.600 165.000 69.900 ;
        RECT 160.100 68.000 160.500 69.500 ;
        RECT 162.200 68.500 162.600 69.500 ;
        RECT 155.800 67.900 157.800 68.000 ;
        RECT 155.100 67.200 155.400 67.900 ;
        RECT 155.900 67.700 157.700 67.900 ;
        RECT 159.700 67.700 160.500 68.000 ;
        RECT 159.700 67.500 160.100 67.700 ;
        RECT 157.000 67.200 157.400 67.400 ;
        RECT 159.700 67.200 160.000 67.500 ;
        RECT 162.300 67.400 162.600 68.500 ;
        RECT 163.000 67.900 163.400 69.600 ;
        RECT 163.800 67.900 164.200 69.300 ;
        RECT 164.600 68.000 165.000 69.600 ;
        RECT 166.200 68.000 166.600 69.900 ;
        RECT 167.800 68.900 168.200 69.900 ;
        RECT 164.600 67.900 166.600 68.000 ;
        RECT 167.000 68.100 167.400 68.200 ;
        RECT 167.800 68.100 168.100 68.900 ;
        RECT 154.200 67.100 154.600 67.200 ;
        RECT 155.000 67.100 156.300 67.200 ;
        RECT 154.200 66.800 156.300 67.100 ;
        RECT 157.000 66.900 157.800 67.200 ;
        RECT 157.400 66.800 157.800 66.900 ;
        RECT 159.000 66.800 160.000 67.200 ;
        RECT 160.500 67.100 162.600 67.400 ;
        RECT 163.800 67.200 164.100 67.900 ;
        RECT 164.700 67.700 166.500 67.900 ;
        RECT 167.000 67.800 168.100 68.100 ;
        RECT 168.600 67.800 169.000 68.600 ;
        RECT 165.800 67.200 166.200 67.400 ;
        RECT 167.800 67.200 168.100 67.800 ;
        RECT 169.400 67.700 169.800 69.900 ;
        RECT 171.500 69.200 172.100 69.900 ;
        RECT 171.500 68.900 172.200 69.200 ;
        RECT 173.800 68.900 174.200 69.900 ;
        RECT 176.000 69.200 176.400 69.900 ;
        RECT 176.000 68.900 177.000 69.200 ;
        RECT 171.800 68.500 172.200 68.900 ;
        RECT 173.900 68.600 174.200 68.900 ;
        RECT 173.900 68.300 175.300 68.600 ;
        RECT 174.900 68.200 175.300 68.300 ;
        RECT 175.800 67.800 176.200 68.600 ;
        RECT 176.600 68.500 177.000 68.900 ;
        RECT 170.900 67.700 171.300 67.800 ;
        RECT 169.400 67.400 171.300 67.700 ;
        RECT 160.500 66.900 161.000 67.100 ;
        RECT 154.200 66.100 154.600 66.200 ;
        RECT 151.800 65.800 152.600 66.100 ;
        RECT 153.400 65.800 154.600 66.100 ;
        RECT 152.200 65.600 152.600 65.800 ;
        RECT 143.100 65.100 144.200 65.200 ;
        RECT 137.100 62.200 138.100 65.100 ;
        RECT 136.600 61.800 138.100 62.200 ;
        RECT 137.100 61.100 138.100 61.800 ;
        RECT 142.700 64.800 144.200 65.100 ;
        RECT 148.900 64.900 150.600 65.200 ;
        RECT 154.200 65.100 154.500 65.800 ;
        RECT 155.000 65.100 155.400 65.200 ;
        RECT 156.000 65.100 156.300 66.800 ;
        RECT 156.600 66.100 157.000 66.600 ;
        RECT 158.200 66.100 158.600 66.200 ;
        RECT 159.000 66.100 159.400 66.200 ;
        RECT 156.600 65.800 159.400 66.100 ;
        RECT 159.000 65.400 159.400 65.800 ;
        RECT 150.200 64.800 150.600 64.900 ;
        RECT 151.800 64.800 153.800 65.100 ;
        RECT 142.700 61.100 143.700 64.800 ;
        RECT 145.500 64.400 147.300 64.700 ;
        RECT 145.500 64.100 145.800 64.400 ;
        RECT 145.400 61.100 145.800 64.100 ;
        RECT 147.000 64.100 147.300 64.400 ;
        RECT 147.900 64.500 149.700 64.600 ;
        RECT 150.200 64.500 150.500 64.800 ;
        RECT 147.900 64.300 149.800 64.500 ;
        RECT 147.900 64.100 148.200 64.300 ;
        RECT 147.000 61.400 147.400 64.100 ;
        RECT 147.800 61.700 148.200 64.100 ;
        RECT 148.600 61.400 149.000 64.000 ;
        RECT 149.400 61.500 149.800 64.300 ;
        RECT 150.200 61.700 150.600 64.500 ;
        RECT 147.000 61.100 149.000 61.400 ;
        RECT 149.500 61.400 149.800 61.500 ;
        RECT 151.000 61.500 151.400 64.500 ;
        RECT 151.000 61.400 151.300 61.500 ;
        RECT 149.500 61.100 151.300 61.400 ;
        RECT 151.800 61.100 152.200 64.800 ;
        RECT 153.400 61.100 153.800 64.800 ;
        RECT 154.200 61.100 154.600 65.100 ;
        RECT 155.000 64.800 155.700 65.100 ;
        RECT 156.000 64.800 156.500 65.100 ;
        RECT 155.400 64.200 155.700 64.800 ;
        RECT 155.400 63.800 155.800 64.200 ;
        RECT 156.100 61.100 156.500 64.800 ;
        RECT 159.700 64.900 160.000 66.800 ;
        RECT 160.300 66.500 161.000 66.900 ;
        RECT 160.700 65.500 161.000 66.500 ;
        RECT 161.400 65.800 161.800 66.600 ;
        RECT 162.200 65.800 162.600 66.600 ;
        RECT 163.000 66.400 163.400 67.200 ;
        RECT 163.800 66.900 165.000 67.200 ;
        RECT 165.800 66.900 166.600 67.200 ;
        RECT 164.600 66.800 165.000 66.900 ;
        RECT 166.200 66.800 166.600 66.900 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 163.800 65.800 164.200 66.600 ;
        RECT 160.700 65.200 162.600 65.500 ;
        RECT 159.700 64.600 160.500 64.900 ;
        RECT 160.100 62.200 160.500 64.600 ;
        RECT 162.300 63.500 162.600 65.200 ;
        RECT 164.700 65.100 165.000 66.800 ;
        RECT 165.400 65.800 165.800 66.600 ;
        RECT 167.000 65.400 167.400 66.200 ;
        RECT 167.800 65.100 168.100 66.800 ;
        RECT 169.400 65.700 169.800 67.400 ;
        RECT 172.900 67.100 173.300 67.200 ;
        RECT 174.200 67.100 174.600 67.200 ;
        RECT 175.800 67.100 176.100 67.800 ;
        RECT 178.200 67.500 178.600 69.900 ;
        RECT 179.000 67.800 179.400 68.600 ;
        RECT 177.400 67.100 178.200 67.200 ;
        RECT 172.700 66.800 178.200 67.100 ;
        RECT 171.800 66.400 172.200 66.500 ;
        RECT 170.300 66.100 172.200 66.400 ;
        RECT 170.300 66.000 170.700 66.100 ;
        RECT 171.100 65.700 171.500 65.800 ;
        RECT 169.400 65.400 171.500 65.700 ;
        RECT 159.800 61.800 160.500 62.200 ;
        RECT 160.100 61.100 160.500 61.800 ;
        RECT 162.200 61.500 162.600 63.500 ;
        RECT 164.300 62.200 165.300 65.100 ;
        RECT 163.800 61.800 165.300 62.200 ;
        RECT 164.300 61.100 165.300 61.800 ;
        RECT 167.300 64.700 168.200 65.100 ;
        RECT 167.300 61.100 167.700 64.700 ;
        RECT 169.400 61.100 169.800 65.400 ;
        RECT 172.700 65.200 173.000 66.800 ;
        RECT 176.300 66.700 176.700 66.800 ;
        RECT 177.100 66.200 177.500 66.300 ;
        RECT 173.400 66.100 173.800 66.200 ;
        RECT 175.000 66.100 177.500 66.200 ;
        RECT 173.400 65.900 177.500 66.100 ;
        RECT 173.400 65.800 175.400 65.900 ;
        RECT 175.800 65.500 178.600 65.600 ;
        RECT 175.700 65.400 178.600 65.500 ;
        RECT 171.800 64.900 173.000 65.200 ;
        RECT 173.700 65.300 178.600 65.400 ;
        RECT 173.700 65.100 176.100 65.300 ;
        RECT 171.800 64.400 172.100 64.900 ;
        RECT 171.400 64.000 172.100 64.400 ;
        RECT 172.900 64.500 173.300 64.600 ;
        RECT 173.700 64.500 174.000 65.100 ;
        RECT 172.900 64.200 174.000 64.500 ;
        RECT 174.300 64.500 177.000 64.800 ;
        RECT 174.300 64.400 174.700 64.500 ;
        RECT 176.600 64.400 177.000 64.500 ;
        RECT 173.500 63.700 173.900 63.800 ;
        RECT 174.900 63.700 175.300 63.800 ;
        RECT 171.800 63.100 172.200 63.500 ;
        RECT 173.500 63.400 175.300 63.700 ;
        RECT 173.900 63.100 174.200 63.400 ;
        RECT 176.600 63.100 177.000 63.500 ;
        RECT 171.500 61.100 172.100 63.100 ;
        RECT 173.800 61.100 174.200 63.100 ;
        RECT 176.000 62.800 177.000 63.100 ;
        RECT 176.000 61.100 176.400 62.800 ;
        RECT 178.200 61.100 178.600 65.300 ;
        RECT 179.800 61.100 180.200 69.900 ;
        RECT 2.500 56.400 2.900 59.900 ;
        RECT 4.600 57.500 5.000 59.500 ;
        RECT 2.100 56.100 2.900 56.400 ;
        RECT 1.400 54.800 1.800 55.600 ;
        RECT 2.100 54.200 2.400 56.100 ;
        RECT 4.700 55.800 5.000 57.500 ;
        RECT 3.100 55.500 5.000 55.800 ;
        RECT 3.100 54.500 3.400 55.500 ;
        RECT 1.400 53.800 2.400 54.200 ;
        RECT 2.700 54.100 3.400 54.500 ;
        RECT 3.800 54.400 4.200 55.200 ;
        RECT 4.600 54.400 5.000 55.200 ;
        RECT 5.400 55.100 5.800 59.900 ;
        RECT 7.000 59.600 9.000 59.900 ;
        RECT 7.000 55.900 7.400 59.600 ;
        RECT 7.800 55.900 8.200 59.300 ;
        RECT 8.600 56.200 9.000 59.600 ;
        RECT 10.200 56.200 10.600 59.900 ;
        RECT 8.600 55.900 10.600 56.200 ;
        RECT 7.900 55.600 8.200 55.900 ;
        RECT 11.000 55.700 11.400 59.900 ;
        RECT 13.200 58.200 13.600 59.900 ;
        RECT 12.600 57.900 13.600 58.200 ;
        RECT 15.400 57.900 15.800 59.900 ;
        RECT 17.500 57.900 18.100 59.900 ;
        RECT 12.600 57.500 13.000 57.900 ;
        RECT 15.400 57.600 15.700 57.900 ;
        RECT 14.300 57.300 16.100 57.600 ;
        RECT 17.400 57.500 17.800 57.900 ;
        RECT 14.300 57.200 14.700 57.300 ;
        RECT 15.700 57.200 16.100 57.300 ;
        RECT 12.600 56.500 13.000 56.600 ;
        RECT 14.900 56.500 15.300 56.600 ;
        RECT 12.600 56.200 15.300 56.500 ;
        RECT 15.600 56.500 16.700 56.800 ;
        RECT 15.600 55.900 15.900 56.500 ;
        RECT 16.300 56.400 16.700 56.500 ;
        RECT 17.500 56.600 18.200 57.000 ;
        RECT 17.500 56.100 17.800 56.600 ;
        RECT 13.500 55.700 15.900 55.900 ;
        RECT 11.000 55.600 15.900 55.700 ;
        RECT 16.600 55.800 17.800 56.100 ;
        RECT 6.200 55.100 6.600 55.200 ;
        RECT 5.400 54.800 6.600 55.100 ;
        RECT 7.000 54.800 7.400 55.600 ;
        RECT 7.900 55.300 8.900 55.600 ;
        RECT 11.000 55.500 13.900 55.600 ;
        RECT 11.000 55.400 13.800 55.500 ;
        RECT 8.600 55.200 8.900 55.300 ;
        RECT 9.800 55.200 10.200 55.400 ;
        RECT 16.600 55.200 16.900 55.800 ;
        RECT 19.800 55.600 20.200 59.900 ;
        RECT 20.600 55.800 21.000 56.600 ;
        RECT 18.100 55.300 20.200 55.600 ;
        RECT 18.100 55.200 18.500 55.300 ;
        RECT 8.600 54.800 9.000 55.200 ;
        RECT 9.800 54.900 10.600 55.200 ;
        RECT 14.200 55.100 14.600 55.200 ;
        RECT 10.200 54.800 10.600 54.900 ;
        RECT 12.100 54.800 14.600 55.100 ;
        RECT 16.600 54.800 17.000 55.200 ;
        RECT 18.900 54.900 19.300 55.000 ;
        RECT 2.100 53.500 2.400 53.800 ;
        RECT 2.900 53.900 3.400 54.100 ;
        RECT 2.900 53.600 5.000 53.900 ;
        RECT 2.100 53.300 2.500 53.500 ;
        RECT 2.100 53.000 2.900 53.300 ;
        RECT 2.500 52.200 2.900 53.000 ;
        RECT 4.700 52.500 5.000 53.600 ;
        RECT 2.500 51.800 3.400 52.200 ;
        RECT 2.500 51.500 2.900 51.800 ;
        RECT 4.600 51.500 5.000 52.500 ;
        RECT 5.400 51.100 5.800 54.800 ;
        RECT 7.900 54.400 8.300 54.800 ;
        RECT 7.900 54.200 8.200 54.400 ;
        RECT 7.800 54.100 8.200 54.200 ;
        RECT 6.200 53.800 8.200 54.100 ;
        RECT 6.200 53.200 6.500 53.800 ;
        RECT 6.200 52.400 6.600 53.200 ;
        RECT 8.600 53.100 8.900 54.800 ;
        RECT 12.100 54.700 12.500 54.800 ;
        RECT 13.400 54.700 13.800 54.800 ;
        RECT 9.400 53.800 9.800 54.600 ;
        RECT 12.900 54.200 13.300 54.300 ;
        RECT 16.600 54.200 16.900 54.800 ;
        RECT 17.400 54.600 19.300 54.900 ;
        RECT 17.400 54.500 17.800 54.600 ;
        RECT 11.400 53.900 16.900 54.200 ;
        RECT 11.400 53.800 12.200 53.900 ;
        RECT 8.300 51.100 9.100 53.100 ;
        RECT 11.000 51.100 11.400 53.500 ;
        RECT 13.500 52.800 13.800 53.900 ;
        RECT 16.300 53.800 16.700 53.900 ;
        RECT 19.800 53.600 20.200 55.300 ;
        RECT 18.300 53.300 20.200 53.600 ;
        RECT 18.300 53.200 18.700 53.300 ;
        RECT 12.600 52.100 13.000 52.500 ;
        RECT 13.400 52.400 13.800 52.800 ;
        RECT 14.300 52.700 14.700 52.800 ;
        RECT 14.300 52.400 15.700 52.700 ;
        RECT 15.400 52.100 15.700 52.400 ;
        RECT 17.400 52.100 17.800 52.500 ;
        RECT 12.600 51.800 13.600 52.100 ;
        RECT 13.200 51.100 13.600 51.800 ;
        RECT 15.400 51.100 15.800 52.100 ;
        RECT 17.400 51.800 18.100 52.100 ;
        RECT 17.500 51.100 18.100 51.800 ;
        RECT 19.800 51.100 20.200 53.300 ;
        RECT 21.400 53.100 21.800 59.900 ;
        RECT 23.000 57.100 23.400 57.200 ;
        RECT 23.800 57.100 24.200 59.900 ;
        RECT 23.000 56.800 24.200 57.100 ;
        RECT 22.200 54.100 22.600 54.200 ;
        RECT 23.000 54.100 23.400 54.200 ;
        RECT 22.200 53.800 23.400 54.100 ;
        RECT 22.200 53.400 22.600 53.800 ;
        RECT 23.000 53.400 23.400 53.800 ;
        RECT 20.900 52.800 21.800 53.100 ;
        RECT 23.800 53.100 24.200 56.800 ;
        RECT 24.600 55.800 25.000 56.600 ;
        RECT 25.400 56.200 25.800 59.900 ;
        RECT 27.000 56.200 27.400 59.900 ;
        RECT 25.400 55.900 27.400 56.200 ;
        RECT 27.800 55.800 28.200 59.900 ;
        RECT 28.900 56.300 29.300 59.900 ;
        RECT 28.900 55.900 29.800 56.300 ;
        RECT 25.800 55.200 26.200 55.400 ;
        RECT 27.800 55.200 28.100 55.800 ;
        RECT 25.400 54.900 26.200 55.200 ;
        RECT 27.000 54.900 28.200 55.200 ;
        RECT 25.400 54.800 25.800 54.900 ;
        RECT 26.200 53.800 26.600 54.600 ;
        RECT 27.000 53.100 27.300 54.900 ;
        RECT 27.800 54.800 28.200 54.900 ;
        RECT 28.600 54.800 29.000 55.600 ;
        RECT 29.400 54.200 29.700 55.900 ;
        RECT 31.000 55.700 31.400 59.900 ;
        RECT 33.200 58.200 33.600 59.900 ;
        RECT 32.600 57.900 33.600 58.200 ;
        RECT 35.400 57.900 35.800 59.900 ;
        RECT 37.500 57.900 38.100 59.900 ;
        RECT 32.600 57.500 33.000 57.900 ;
        RECT 35.400 57.600 35.700 57.900 ;
        RECT 34.300 57.300 36.100 57.600 ;
        RECT 37.400 57.500 37.800 57.900 ;
        RECT 34.300 57.200 34.700 57.300 ;
        RECT 35.700 57.200 36.100 57.300 ;
        RECT 39.800 57.100 40.200 59.900 ;
        RECT 40.600 57.100 41.000 57.200 ;
        RECT 32.600 56.500 33.000 56.600 ;
        RECT 34.900 56.500 35.300 56.600 ;
        RECT 32.600 56.200 35.300 56.500 ;
        RECT 35.600 56.500 36.700 56.800 ;
        RECT 35.600 55.900 35.900 56.500 ;
        RECT 36.300 56.400 36.700 56.500 ;
        RECT 37.500 56.600 38.200 57.000 ;
        RECT 39.800 56.800 41.000 57.100 ;
        RECT 37.500 56.100 37.800 56.600 ;
        RECT 33.500 55.700 35.900 55.900 ;
        RECT 31.000 55.600 35.900 55.700 ;
        RECT 36.600 55.800 37.800 56.100 ;
        RECT 31.000 55.500 33.900 55.600 ;
        RECT 31.000 55.400 33.800 55.500 ;
        RECT 34.200 55.100 34.600 55.200 ;
        RECT 32.100 54.800 34.600 55.100 ;
        RECT 32.100 54.700 32.500 54.800 ;
        RECT 33.400 54.700 33.800 54.800 ;
        RECT 32.900 54.200 33.300 54.300 ;
        RECT 36.600 54.200 36.900 55.800 ;
        RECT 39.800 55.600 40.200 56.800 ;
        RECT 42.200 56.200 42.600 59.900 ;
        RECT 43.800 59.600 45.800 59.900 ;
        RECT 43.800 56.200 44.200 59.600 ;
        RECT 42.200 55.900 44.200 56.200 ;
        RECT 44.600 55.900 45.000 59.300 ;
        RECT 45.400 55.900 45.800 59.600 ;
        RECT 46.200 57.900 46.600 59.900 ;
        RECT 46.300 57.800 46.600 57.900 ;
        RECT 47.800 57.900 48.200 59.900 ;
        RECT 47.800 57.800 48.100 57.900 ;
        RECT 46.300 57.500 48.100 57.800 ;
        RECT 46.300 56.200 46.600 57.500 ;
        RECT 47.000 56.400 47.400 57.200 ;
        RECT 44.600 55.600 44.900 55.900 ;
        RECT 46.200 55.800 46.600 56.200 ;
        RECT 38.100 55.300 40.200 55.600 ;
        RECT 38.100 55.200 38.500 55.300 ;
        RECT 38.900 54.900 39.300 55.000 ;
        RECT 37.400 54.600 39.300 54.900 ;
        RECT 37.400 54.500 37.800 54.600 ;
        RECT 29.400 53.800 29.800 54.200 ;
        RECT 31.400 53.900 37.000 54.200 ;
        RECT 31.400 53.800 32.200 53.900 ;
        RECT 27.800 53.100 28.200 53.200 ;
        RECT 29.400 53.100 29.700 53.800 ;
        RECT 23.800 52.800 24.700 53.100 ;
        RECT 20.900 52.200 21.300 52.800 ;
        RECT 20.600 51.800 21.300 52.200 ;
        RECT 20.900 51.100 21.300 51.800 ;
        RECT 24.300 51.100 24.700 52.800 ;
        RECT 27.000 51.100 27.400 53.100 ;
        RECT 27.800 52.800 29.700 53.100 ;
        RECT 27.700 52.400 28.100 52.800 ;
        RECT 29.400 52.100 29.700 52.800 ;
        RECT 30.200 52.400 30.600 53.200 ;
        RECT 29.400 51.100 29.800 52.100 ;
        RECT 31.000 51.100 31.400 53.500 ;
        RECT 33.500 52.800 33.800 53.900 ;
        RECT 36.300 53.800 37.000 53.900 ;
        RECT 39.800 53.600 40.200 55.300 ;
        RECT 42.600 55.200 43.000 55.400 ;
        RECT 43.900 55.300 44.900 55.600 ;
        RECT 43.900 55.200 44.200 55.300 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 42.200 55.100 43.000 55.200 ;
        RECT 40.600 54.900 43.000 55.100 ;
        RECT 40.600 54.800 42.600 54.900 ;
        RECT 43.800 54.800 44.200 55.200 ;
        RECT 45.400 54.800 45.800 55.600 ;
        RECT 43.000 53.800 43.400 54.600 ;
        RECT 38.300 53.300 40.200 53.600 ;
        RECT 38.300 53.200 38.700 53.300 ;
        RECT 32.600 52.100 33.000 52.500 ;
        RECT 33.400 52.400 33.800 52.800 ;
        RECT 34.300 52.700 34.700 52.800 ;
        RECT 34.300 52.400 35.700 52.700 ;
        RECT 35.400 52.100 35.700 52.400 ;
        RECT 37.400 52.100 37.800 52.500 ;
        RECT 32.600 51.800 33.600 52.100 ;
        RECT 33.200 51.100 33.600 51.800 ;
        RECT 35.400 51.100 35.800 52.100 ;
        RECT 37.400 51.800 38.100 52.100 ;
        RECT 37.500 51.100 38.100 51.800 ;
        RECT 39.800 51.100 40.200 53.300 ;
        RECT 43.900 53.100 44.200 54.800 ;
        RECT 44.500 54.400 44.900 54.800 ;
        RECT 44.600 54.200 44.900 54.400 ;
        RECT 46.300 54.200 46.600 55.800 ;
        RECT 48.600 55.400 49.000 56.200 ;
        RECT 49.400 55.800 49.800 56.600 ;
        RECT 47.400 54.800 48.200 55.200 ;
        RECT 50.200 55.100 50.600 59.900 ;
        RECT 49.400 54.800 50.600 55.100 ;
        RECT 49.400 54.200 49.700 54.800 ;
        RECT 44.600 53.800 45.000 54.200 ;
        RECT 46.300 54.100 47.100 54.200 ;
        RECT 46.300 53.900 47.200 54.100 ;
        RECT 43.700 51.100 44.500 53.100 ;
        RECT 46.800 51.100 47.200 53.900 ;
        RECT 49.400 53.800 49.800 54.200 ;
        RECT 50.200 53.100 50.600 54.800 ;
        RECT 51.000 54.100 51.400 54.200 ;
        RECT 51.800 54.100 52.200 54.200 ;
        RECT 51.000 53.800 52.200 54.100 ;
        RECT 51.000 53.400 51.400 53.800 ;
        RECT 49.700 52.800 50.600 53.100 ;
        RECT 49.700 51.100 50.100 52.800 ;
        RECT 52.600 51.100 53.000 59.900 ;
        RECT 55.500 56.300 55.900 59.900 ;
        RECT 55.000 55.900 55.900 56.300 ;
        RECT 55.100 54.200 55.400 55.900 ;
        RECT 56.600 55.600 57.000 59.900 ;
        RECT 58.700 57.900 59.300 59.900 ;
        RECT 61.000 57.900 61.400 59.900 ;
        RECT 63.200 58.200 63.600 59.900 ;
        RECT 63.200 57.900 64.200 58.200 ;
        RECT 59.000 57.500 59.400 57.900 ;
        RECT 61.100 57.600 61.400 57.900 ;
        RECT 60.700 57.300 62.500 57.600 ;
        RECT 63.800 57.500 64.200 57.900 ;
        RECT 60.700 57.200 61.100 57.300 ;
        RECT 62.100 57.200 62.500 57.300 ;
        RECT 58.600 56.600 59.300 57.000 ;
        RECT 59.000 56.100 59.300 56.600 ;
        RECT 60.100 56.500 61.200 56.800 ;
        RECT 60.100 56.400 60.500 56.500 ;
        RECT 59.000 55.800 60.200 56.100 ;
        RECT 55.800 54.800 56.200 55.600 ;
        RECT 56.600 55.300 58.700 55.600 ;
        RECT 53.400 53.400 53.800 54.200 ;
        RECT 55.000 53.800 55.400 54.200 ;
        RECT 54.200 52.400 54.600 53.200 ;
        RECT 55.100 52.200 55.400 53.800 ;
        RECT 55.000 51.100 55.400 52.200 ;
        RECT 56.600 53.600 57.000 55.300 ;
        RECT 58.300 55.200 58.700 55.300 ;
        RECT 57.500 54.900 57.900 55.000 ;
        RECT 57.500 54.600 59.400 54.900 ;
        RECT 59.000 54.500 59.400 54.600 ;
        RECT 59.900 54.200 60.200 55.800 ;
        RECT 60.900 55.900 61.200 56.500 ;
        RECT 61.500 56.500 61.900 56.600 ;
        RECT 63.800 56.500 64.200 56.600 ;
        RECT 61.500 56.200 64.200 56.500 ;
        RECT 60.900 55.700 63.300 55.900 ;
        RECT 65.400 55.700 65.800 59.900 ;
        RECT 66.500 59.200 66.900 59.900 ;
        RECT 66.200 58.800 66.900 59.200 ;
        RECT 66.500 56.300 66.900 58.800 ;
        RECT 69.900 56.300 70.300 59.900 ;
        RECT 66.500 55.900 67.400 56.300 ;
        RECT 69.400 55.900 70.300 56.300 ;
        RECT 71.300 59.200 71.700 59.900 ;
        RECT 71.300 58.800 72.200 59.200 ;
        RECT 71.300 56.300 71.700 58.800 ;
        RECT 73.400 57.500 73.800 59.500 ;
        RECT 71.300 55.900 72.200 56.300 ;
        RECT 60.900 55.600 65.800 55.700 ;
        RECT 62.900 55.500 65.800 55.600 ;
        RECT 63.000 55.400 65.800 55.500 ;
        RECT 62.200 55.100 62.600 55.200 ;
        RECT 62.200 54.800 64.700 55.100 ;
        RECT 66.200 54.800 66.600 55.600 ;
        RECT 64.300 54.700 64.700 54.800 ;
        RECT 63.500 54.200 63.900 54.300 ;
        RECT 67.000 54.200 67.300 55.900 ;
        RECT 69.500 54.200 69.800 55.900 ;
        RECT 70.200 55.100 70.600 55.600 ;
        RECT 71.000 55.100 71.400 55.600 ;
        RECT 70.200 54.800 71.400 55.100 ;
        RECT 59.900 53.900 65.400 54.200 ;
        RECT 60.100 53.800 60.500 53.900 ;
        RECT 61.400 53.800 61.800 53.900 ;
        RECT 56.600 53.300 58.500 53.600 ;
        RECT 56.600 51.100 57.000 53.300 ;
        RECT 58.100 53.200 58.500 53.300 ;
        RECT 63.000 52.800 63.300 53.900 ;
        RECT 64.600 53.800 65.400 53.900 ;
        RECT 67.000 53.800 67.400 54.200 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 69.400 54.100 69.800 54.200 ;
        RECT 68.600 53.800 69.800 54.100 ;
        RECT 62.100 52.700 62.500 52.800 ;
        RECT 59.000 52.100 59.400 52.500 ;
        RECT 61.100 52.400 62.500 52.700 ;
        RECT 63.000 52.400 63.400 52.800 ;
        RECT 61.100 52.100 61.400 52.400 ;
        RECT 63.800 52.100 64.200 52.500 ;
        RECT 58.700 51.800 59.400 52.100 ;
        RECT 58.700 51.100 59.300 51.800 ;
        RECT 61.000 51.100 61.400 52.100 ;
        RECT 63.200 51.800 64.200 52.100 ;
        RECT 63.200 51.100 63.600 51.800 ;
        RECT 65.400 51.100 65.800 53.500 ;
        RECT 67.000 52.100 67.300 53.800 ;
        RECT 67.800 52.400 68.200 53.200 ;
        RECT 68.600 52.400 69.000 53.200 ;
        RECT 69.500 52.100 69.800 53.800 ;
        RECT 67.000 51.100 67.400 52.100 ;
        RECT 69.400 51.100 69.800 52.100 ;
        RECT 71.800 54.200 72.100 55.900 ;
        RECT 73.400 55.800 73.700 57.500 ;
        RECT 75.500 56.400 75.900 59.900 ;
        RECT 75.500 56.100 76.300 56.400 ;
        RECT 73.400 55.500 75.300 55.800 ;
        RECT 73.400 54.400 73.800 55.200 ;
        RECT 74.200 54.400 74.600 55.200 ;
        RECT 75.000 54.500 75.300 55.500 ;
        RECT 71.800 53.800 72.200 54.200 ;
        RECT 75.000 54.100 75.700 54.500 ;
        RECT 76.000 54.200 76.300 56.100 ;
        RECT 76.600 55.100 77.000 55.600 ;
        RECT 78.200 55.100 78.600 59.900 ;
        RECT 79.800 56.200 80.200 59.900 ;
        RECT 81.400 59.600 83.400 59.900 ;
        RECT 81.400 56.200 81.800 59.600 ;
        RECT 79.800 55.900 81.800 56.200 ;
        RECT 82.200 55.900 82.600 59.300 ;
        RECT 83.000 55.900 83.400 59.600 ;
        RECT 82.200 55.600 82.500 55.900 ;
        RECT 83.800 55.600 84.200 59.900 ;
        RECT 85.900 57.900 86.500 59.900 ;
        RECT 88.200 57.900 88.600 59.900 ;
        RECT 90.400 58.200 90.800 59.900 ;
        RECT 90.400 57.900 91.400 58.200 ;
        RECT 86.200 57.500 86.600 57.900 ;
        RECT 88.300 57.600 88.600 57.900 ;
        RECT 87.900 57.300 89.700 57.600 ;
        RECT 91.000 57.500 91.400 57.900 ;
        RECT 87.900 57.200 88.300 57.300 ;
        RECT 89.300 57.200 89.700 57.300 ;
        RECT 85.800 56.600 86.500 57.000 ;
        RECT 86.200 56.100 86.500 56.600 ;
        RECT 87.300 56.500 88.400 56.800 ;
        RECT 87.300 56.400 87.700 56.500 ;
        RECT 86.200 55.800 87.400 56.100 ;
        RECT 80.200 55.200 80.600 55.400 ;
        RECT 81.500 55.300 82.500 55.600 ;
        RECT 81.500 55.200 81.800 55.300 ;
        RECT 76.600 54.800 78.600 55.100 ;
        RECT 79.000 55.100 79.400 55.200 ;
        RECT 79.800 55.100 80.600 55.200 ;
        RECT 79.000 54.900 80.600 55.100 ;
        RECT 79.000 54.800 80.200 54.900 ;
        RECT 81.400 54.800 81.800 55.200 ;
        RECT 83.000 54.800 83.400 55.600 ;
        RECT 83.800 55.300 85.900 55.600 ;
        RECT 75.000 53.900 75.500 54.100 ;
        RECT 71.800 52.100 72.100 53.800 ;
        RECT 73.400 53.600 75.500 53.900 ;
        RECT 76.000 53.800 77.000 54.200 ;
        RECT 72.600 52.400 73.000 53.200 ;
        RECT 73.400 52.500 73.700 53.600 ;
        RECT 76.000 53.500 76.300 53.800 ;
        RECT 75.900 53.300 76.300 53.500 ;
        RECT 75.500 53.000 76.300 53.300 ;
        RECT 71.800 51.100 72.200 52.100 ;
        RECT 73.400 51.500 73.800 52.500 ;
        RECT 75.500 52.200 75.900 53.000 ;
        RECT 75.000 51.800 75.900 52.200 ;
        RECT 75.500 51.500 75.900 51.800 ;
        RECT 78.200 51.100 78.600 54.800 ;
        RECT 79.800 54.100 80.200 54.200 ;
        RECT 80.600 54.100 81.000 54.600 ;
        RECT 79.000 53.800 81.000 54.100 ;
        RECT 79.000 53.200 79.300 53.800 ;
        RECT 79.000 52.400 79.400 53.200 ;
        RECT 81.500 53.100 81.800 54.800 ;
        RECT 82.100 54.400 82.500 54.800 ;
        RECT 82.200 54.200 82.500 54.400 ;
        RECT 82.200 53.800 82.600 54.200 ;
        RECT 83.800 53.600 84.200 55.300 ;
        RECT 85.500 55.200 85.900 55.300 ;
        RECT 84.700 54.900 85.100 55.000 ;
        RECT 84.700 54.600 86.600 54.900 ;
        RECT 86.200 54.500 86.600 54.600 ;
        RECT 87.100 54.200 87.400 55.800 ;
        RECT 88.100 55.900 88.400 56.500 ;
        RECT 88.700 56.500 89.100 56.600 ;
        RECT 91.000 56.500 91.400 56.600 ;
        RECT 88.700 56.200 91.400 56.500 ;
        RECT 88.100 55.700 90.500 55.900 ;
        RECT 92.600 55.700 93.000 59.900 ;
        RECT 95.000 56.200 95.400 59.900 ;
        RECT 96.600 56.200 97.000 59.900 ;
        RECT 95.000 55.900 97.000 56.200 ;
        RECT 97.400 55.900 97.800 59.900 ;
        RECT 99.500 56.300 99.900 59.900 ;
        RECT 99.000 55.900 99.900 56.300 ;
        RECT 88.100 55.600 93.000 55.700 ;
        RECT 90.100 55.500 93.000 55.600 ;
        RECT 90.200 55.400 93.000 55.500 ;
        RECT 95.400 55.200 95.800 55.400 ;
        RECT 97.400 55.200 97.700 55.900 ;
        RECT 89.400 55.100 89.800 55.200 ;
        RECT 89.400 54.800 91.900 55.100 ;
        RECT 95.000 54.900 95.800 55.200 ;
        RECT 96.600 54.900 97.800 55.200 ;
        RECT 95.000 54.800 95.400 54.900 ;
        RECT 90.200 54.700 90.600 54.800 ;
        RECT 91.500 54.700 91.900 54.800 ;
        RECT 90.700 54.200 91.100 54.300 ;
        RECT 87.100 53.900 92.600 54.200 ;
        RECT 87.300 53.800 87.700 53.900 ;
        RECT 88.600 53.800 89.000 53.900 ;
        RECT 83.800 53.300 85.700 53.600 ;
        RECT 81.300 51.100 82.100 53.100 ;
        RECT 83.800 51.100 84.200 53.300 ;
        RECT 85.300 53.200 85.700 53.300 ;
        RECT 90.200 52.800 90.500 53.900 ;
        RECT 91.800 53.800 92.600 53.900 ;
        RECT 95.800 53.800 96.200 54.600 ;
        RECT 89.300 52.700 89.700 52.800 ;
        RECT 86.200 52.100 86.600 52.500 ;
        RECT 88.300 52.400 89.700 52.700 ;
        RECT 90.200 52.400 90.600 52.800 ;
        RECT 88.300 52.100 88.600 52.400 ;
        RECT 91.000 52.100 91.400 52.500 ;
        RECT 85.900 51.800 86.600 52.100 ;
        RECT 85.900 51.100 86.500 51.800 ;
        RECT 88.200 51.100 88.600 52.100 ;
        RECT 90.400 51.800 91.400 52.100 ;
        RECT 90.400 51.100 90.800 51.800 ;
        RECT 92.600 51.100 93.000 53.500 ;
        RECT 96.600 53.200 96.900 54.900 ;
        RECT 97.400 54.800 97.800 54.900 ;
        RECT 99.100 54.200 99.400 55.900 ;
        RECT 100.600 55.600 101.000 59.900 ;
        RECT 102.700 57.900 103.300 59.900 ;
        RECT 105.000 57.900 105.400 59.900 ;
        RECT 107.200 58.200 107.600 59.900 ;
        RECT 107.200 57.900 108.200 58.200 ;
        RECT 103.000 57.500 103.400 57.900 ;
        RECT 105.100 57.600 105.400 57.900 ;
        RECT 104.700 57.300 106.500 57.600 ;
        RECT 107.800 57.500 108.200 57.900 ;
        RECT 104.700 57.200 105.100 57.300 ;
        RECT 106.100 57.200 106.500 57.300 ;
        RECT 102.600 56.600 103.300 57.000 ;
        RECT 103.000 56.100 103.300 56.600 ;
        RECT 104.100 56.500 105.200 56.800 ;
        RECT 104.100 56.400 104.500 56.500 ;
        RECT 103.000 55.800 104.200 56.100 ;
        RECT 99.800 54.800 100.200 55.600 ;
        RECT 100.600 55.300 102.700 55.600 ;
        RECT 99.000 54.100 99.400 54.200 ;
        RECT 97.400 53.800 99.400 54.100 ;
        RECT 97.400 53.200 97.700 53.800 ;
        RECT 96.600 51.100 97.000 53.200 ;
        RECT 97.400 52.800 97.800 53.200 ;
        RECT 97.300 52.400 97.700 52.800 ;
        RECT 98.200 52.400 98.600 53.200 ;
        RECT 99.100 52.100 99.400 53.800 ;
        RECT 99.000 51.100 99.400 52.100 ;
        RECT 100.600 53.600 101.000 55.300 ;
        RECT 102.300 55.200 102.700 55.300 ;
        RECT 101.500 54.900 101.900 55.000 ;
        RECT 101.500 54.600 103.400 54.900 ;
        RECT 103.000 54.500 103.400 54.600 ;
        RECT 103.900 54.200 104.200 55.800 ;
        RECT 104.900 55.900 105.200 56.500 ;
        RECT 105.500 56.500 105.900 56.600 ;
        RECT 107.800 56.500 108.200 56.600 ;
        RECT 105.500 56.200 108.200 56.500 ;
        RECT 104.900 55.700 107.300 55.900 ;
        RECT 109.400 55.700 109.800 59.900 ;
        RECT 104.900 55.600 109.800 55.700 ;
        RECT 106.900 55.500 109.800 55.600 ;
        RECT 107.000 55.400 109.800 55.500 ;
        RECT 106.200 55.100 106.600 55.200 ;
        RECT 111.000 55.100 111.400 59.900 ;
        RECT 113.700 56.400 114.100 59.900 ;
        RECT 115.800 57.500 116.200 59.500 ;
        RECT 113.300 56.100 114.100 56.400 ;
        RECT 112.600 55.100 113.000 55.600 ;
        RECT 106.200 54.800 108.700 55.100 ;
        RECT 107.000 54.700 107.400 54.800 ;
        RECT 108.300 54.700 108.700 54.800 ;
        RECT 111.000 54.800 113.000 55.100 ;
        RECT 107.500 54.200 107.900 54.300 ;
        RECT 103.900 53.900 109.400 54.200 ;
        RECT 104.100 53.800 104.500 53.900 ;
        RECT 105.400 53.800 105.800 53.900 ;
        RECT 100.600 53.300 102.500 53.600 ;
        RECT 100.600 51.100 101.000 53.300 ;
        RECT 102.100 53.200 102.500 53.300 ;
        RECT 107.000 52.800 107.300 53.900 ;
        RECT 108.600 53.800 109.400 53.900 ;
        RECT 106.100 52.700 106.500 52.800 ;
        RECT 103.000 52.100 103.400 52.500 ;
        RECT 105.100 52.400 106.500 52.700 ;
        RECT 107.000 52.400 107.400 52.800 ;
        RECT 105.100 52.100 105.400 52.400 ;
        RECT 107.800 52.100 108.200 52.500 ;
        RECT 102.700 51.800 103.400 52.100 ;
        RECT 102.700 51.100 103.300 51.800 ;
        RECT 105.000 51.100 105.400 52.100 ;
        RECT 107.200 51.800 108.200 52.100 ;
        RECT 107.200 51.100 107.600 51.800 ;
        RECT 109.400 51.100 109.800 53.500 ;
        RECT 110.200 52.400 110.600 53.200 ;
        RECT 111.000 51.100 111.400 54.800 ;
        RECT 113.300 54.200 113.600 56.100 ;
        RECT 115.900 55.800 116.200 57.500 ;
        RECT 114.300 55.500 116.200 55.800 ;
        RECT 114.300 54.500 114.600 55.500 ;
        RECT 111.800 54.100 112.200 54.200 ;
        RECT 112.600 54.100 113.600 54.200 ;
        RECT 113.900 54.100 114.600 54.500 ;
        RECT 115.000 54.400 115.400 55.200 ;
        RECT 115.800 54.400 116.200 55.200 ;
        RECT 111.800 53.800 113.600 54.100 ;
        RECT 113.300 53.500 113.600 53.800 ;
        RECT 114.100 53.900 114.600 54.100 ;
        RECT 114.100 53.600 116.200 53.900 ;
        RECT 113.300 53.300 113.700 53.500 ;
        RECT 113.300 53.000 114.100 53.300 ;
        RECT 113.700 51.500 114.100 53.000 ;
        RECT 115.900 52.500 116.200 53.600 ;
        RECT 115.800 51.500 116.200 52.500 ;
        RECT 116.600 52.400 117.000 53.200 ;
        RECT 117.400 51.100 117.800 59.900 ;
        RECT 118.200 53.400 118.600 54.200 ;
        RECT 119.000 51.100 119.400 59.900 ;
        RECT 120.700 59.600 122.500 59.900 ;
        RECT 120.700 59.500 121.000 59.600 ;
        RECT 120.600 56.500 121.000 59.500 ;
        RECT 122.200 59.500 122.500 59.600 ;
        RECT 123.000 59.600 125.000 59.900 ;
        RECT 121.400 56.500 121.800 59.300 ;
        RECT 122.200 56.700 122.600 59.500 ;
        RECT 123.000 57.000 123.400 59.600 ;
        RECT 123.800 56.900 124.200 59.300 ;
        RECT 124.600 56.900 125.000 59.600 ;
        RECT 123.800 56.700 124.100 56.900 ;
        RECT 122.200 56.500 124.100 56.700 ;
        RECT 121.500 56.200 121.800 56.500 ;
        RECT 122.300 56.400 124.100 56.500 ;
        RECT 124.700 56.600 125.000 56.900 ;
        RECT 126.200 56.900 126.600 59.900 ;
        RECT 126.200 56.600 126.500 56.900 ;
        RECT 124.700 56.300 126.500 56.600 ;
        RECT 121.400 56.100 121.800 56.200 ;
        RECT 121.400 55.800 123.100 56.100 ;
        RECT 122.800 52.500 123.100 55.800 ;
        RECT 127.000 55.600 127.400 59.900 ;
        RECT 129.100 57.900 129.700 59.900 ;
        RECT 131.400 57.900 131.800 59.900 ;
        RECT 133.600 58.200 134.000 59.900 ;
        RECT 133.600 57.900 134.600 58.200 ;
        RECT 129.400 57.500 129.800 57.900 ;
        RECT 131.500 57.600 131.800 57.900 ;
        RECT 131.100 57.300 132.900 57.600 ;
        RECT 134.200 57.500 134.600 57.900 ;
        RECT 131.100 57.200 131.500 57.300 ;
        RECT 132.500 57.200 132.900 57.300 ;
        RECT 129.000 56.600 129.700 57.000 ;
        RECT 129.400 56.100 129.700 56.600 ;
        RECT 130.500 56.500 131.600 56.800 ;
        RECT 130.500 56.400 130.900 56.500 ;
        RECT 129.400 55.800 130.600 56.100 ;
        RECT 127.000 55.300 129.100 55.600 ;
        RECT 123.400 54.800 124.200 55.200 ;
        RECT 124.200 53.800 125.000 54.200 ;
        RECT 127.000 53.600 127.400 55.300 ;
        RECT 128.700 55.200 129.100 55.300 ;
        RECT 127.900 54.900 128.300 55.000 ;
        RECT 127.900 54.600 129.800 54.900 ;
        RECT 129.400 54.500 129.800 54.600 ;
        RECT 130.300 54.200 130.600 55.800 ;
        RECT 131.300 55.900 131.600 56.500 ;
        RECT 131.900 56.500 132.300 56.600 ;
        RECT 134.200 56.500 134.600 56.600 ;
        RECT 131.900 56.200 134.600 56.500 ;
        RECT 131.300 55.700 133.700 55.900 ;
        RECT 135.800 55.700 136.200 59.900 ;
        RECT 131.300 55.600 136.200 55.700 ;
        RECT 133.300 55.500 136.200 55.600 ;
        RECT 133.400 55.400 136.200 55.500 ;
        RECT 137.400 56.100 137.800 59.900 ;
        RECT 141.700 56.400 142.100 59.900 ;
        RECT 143.800 57.500 144.200 59.500 ;
        RECT 138.200 56.100 138.600 56.200 ;
        RECT 137.400 55.800 138.600 56.100 ;
        RECT 141.300 56.100 142.100 56.400 ;
        RECT 132.600 55.100 133.000 55.200 ;
        RECT 132.600 54.800 135.100 55.100 ;
        RECT 133.400 54.700 133.800 54.800 ;
        RECT 134.700 54.700 135.100 54.800 ;
        RECT 133.900 54.200 134.300 54.300 ;
        RECT 130.300 53.900 135.800 54.200 ;
        RECT 130.500 53.800 130.900 53.900 ;
        RECT 127.000 53.300 128.900 53.600 ;
        RECT 124.900 53.100 125.800 53.200 ;
        RECT 126.200 53.100 126.600 53.200 ;
        RECT 124.900 52.800 126.600 53.100 ;
        RECT 122.800 52.200 124.800 52.500 ;
        RECT 122.800 52.100 123.400 52.200 ;
        RECT 123.000 51.100 123.400 52.100 ;
        RECT 124.500 52.100 124.800 52.200 ;
        RECT 124.500 51.800 125.000 52.100 ;
        RECT 124.600 51.100 125.000 51.800 ;
        RECT 127.000 51.100 127.400 53.300 ;
        RECT 128.500 53.200 128.900 53.300 ;
        RECT 133.400 52.800 133.700 53.900 ;
        RECT 135.000 53.800 135.800 53.900 ;
        RECT 132.500 52.700 132.900 52.800 ;
        RECT 129.400 52.100 129.800 52.500 ;
        RECT 131.500 52.400 132.900 52.700 ;
        RECT 133.400 52.400 133.800 52.800 ;
        RECT 131.500 52.100 131.800 52.400 ;
        RECT 134.200 52.100 134.600 52.500 ;
        RECT 129.100 51.800 129.800 52.100 ;
        RECT 129.100 51.100 129.700 51.800 ;
        RECT 131.400 51.100 131.800 52.100 ;
        RECT 133.600 51.800 134.600 52.100 ;
        RECT 133.600 51.100 134.000 51.800 ;
        RECT 135.800 51.100 136.200 53.500 ;
        RECT 136.600 52.400 137.000 53.200 ;
        RECT 137.400 51.100 137.800 55.800 ;
        RECT 140.600 54.800 141.000 55.600 ;
        RECT 141.300 54.200 141.600 56.100 ;
        RECT 143.900 55.800 144.200 57.500 ;
        RECT 142.300 55.500 144.200 55.800 ;
        RECT 144.600 55.700 145.000 59.900 ;
        RECT 146.800 58.200 147.200 59.900 ;
        RECT 146.200 57.900 147.200 58.200 ;
        RECT 149.000 57.900 149.400 59.900 ;
        RECT 151.100 57.900 151.700 59.900 ;
        RECT 146.200 57.500 146.600 57.900 ;
        RECT 149.000 57.600 149.300 57.900 ;
        RECT 147.900 57.300 149.700 57.600 ;
        RECT 151.000 57.500 151.400 57.900 ;
        RECT 147.900 57.200 148.300 57.300 ;
        RECT 149.300 57.200 149.700 57.300 ;
        RECT 146.200 56.500 146.600 56.600 ;
        RECT 148.500 56.500 148.900 56.600 ;
        RECT 146.200 56.200 148.900 56.500 ;
        RECT 149.200 56.500 150.300 56.800 ;
        RECT 149.200 55.900 149.500 56.500 ;
        RECT 149.900 56.400 150.300 56.500 ;
        RECT 151.100 56.600 151.800 57.000 ;
        RECT 151.100 56.100 151.400 56.600 ;
        RECT 147.100 55.700 149.500 55.900 ;
        RECT 144.600 55.600 149.500 55.700 ;
        RECT 150.200 55.800 151.400 56.100 ;
        RECT 144.600 55.500 147.500 55.600 ;
        RECT 142.300 54.500 142.600 55.500 ;
        RECT 144.600 55.400 147.400 55.500 ;
        RECT 138.200 54.100 138.600 54.200 ;
        RECT 140.600 54.100 141.600 54.200 ;
        RECT 141.900 54.100 142.600 54.500 ;
        RECT 143.000 54.400 143.400 55.200 ;
        RECT 143.800 54.400 144.200 55.200 ;
        RECT 147.800 55.100 148.200 55.200 ;
        RECT 145.700 54.800 148.200 55.100 ;
        RECT 145.700 54.700 146.100 54.800 ;
        RECT 146.500 54.200 146.900 54.300 ;
        RECT 150.200 54.200 150.500 55.800 ;
        RECT 153.400 55.600 153.800 59.900 ;
        RECT 151.700 55.300 153.800 55.600 ;
        RECT 154.200 57.500 154.600 59.500 ;
        RECT 154.200 55.800 154.500 57.500 ;
        RECT 156.300 56.400 156.700 59.900 ;
        RECT 159.000 56.900 159.400 59.900 ;
        RECT 159.100 56.600 159.400 56.900 ;
        RECT 160.600 59.600 162.600 59.900 ;
        RECT 160.600 56.900 161.000 59.600 ;
        RECT 161.400 56.900 161.800 59.300 ;
        RECT 162.200 57.000 162.600 59.600 ;
        RECT 163.100 59.600 164.900 59.900 ;
        RECT 163.100 59.500 163.400 59.600 ;
        RECT 160.600 56.600 160.900 56.900 ;
        RECT 156.300 56.100 157.100 56.400 ;
        RECT 159.100 56.300 160.900 56.600 ;
        RECT 161.500 56.700 161.800 56.900 ;
        RECT 163.000 56.700 163.400 59.500 ;
        RECT 164.600 59.500 164.900 59.600 ;
        RECT 161.500 56.500 163.400 56.700 ;
        RECT 163.800 56.500 164.200 59.300 ;
        RECT 164.600 56.500 165.000 59.500 ;
        RECT 165.400 57.500 165.800 59.500 ;
        RECT 167.500 59.200 167.900 59.900 ;
        RECT 167.500 58.800 168.200 59.200 ;
        RECT 161.500 56.400 163.300 56.500 ;
        RECT 163.800 56.200 164.100 56.500 ;
        RECT 163.800 56.100 164.200 56.200 ;
        RECT 154.200 55.500 156.100 55.800 ;
        RECT 151.700 55.200 152.100 55.300 ;
        RECT 152.500 54.900 152.900 55.000 ;
        RECT 151.000 54.600 152.900 54.900 ;
        RECT 151.000 54.500 151.400 54.600 ;
        RECT 138.200 53.800 141.600 54.100 ;
        RECT 141.300 53.500 141.600 53.800 ;
        RECT 142.100 53.900 142.600 54.100 ;
        RECT 145.000 53.900 150.600 54.200 ;
        RECT 142.100 53.600 144.200 53.900 ;
        RECT 145.000 53.800 145.800 53.900 ;
        RECT 141.300 53.300 141.700 53.500 ;
        RECT 141.300 53.000 142.100 53.300 ;
        RECT 141.700 51.500 142.100 53.000 ;
        RECT 143.900 52.500 144.200 53.600 ;
        RECT 143.800 51.500 144.200 52.500 ;
        RECT 144.600 51.100 145.000 53.500 ;
        RECT 147.100 52.800 147.400 53.900 ;
        RECT 149.900 53.800 150.600 53.900 ;
        RECT 153.400 53.600 153.800 55.300 ;
        RECT 154.200 54.400 154.600 55.200 ;
        RECT 155.000 54.400 155.400 55.200 ;
        RECT 155.800 54.500 156.100 55.500 ;
        RECT 155.800 54.100 156.500 54.500 ;
        RECT 156.800 54.200 157.100 56.100 ;
        RECT 162.500 55.800 164.200 56.100 ;
        RECT 165.400 55.800 165.700 57.500 ;
        RECT 167.500 56.400 167.900 58.800 ;
        RECT 167.500 56.100 168.300 56.400 ;
        RECT 162.500 55.700 163.400 55.800 ;
        RECT 157.400 54.800 157.800 55.600 ;
        RECT 161.400 54.800 162.200 55.200 ;
        RECT 155.800 53.900 156.300 54.100 ;
        RECT 151.900 53.300 153.800 53.600 ;
        RECT 151.900 53.200 152.300 53.300 ;
        RECT 146.200 52.100 146.600 52.500 ;
        RECT 147.000 52.400 147.400 52.800 ;
        RECT 147.900 52.700 148.300 52.800 ;
        RECT 147.900 52.400 149.300 52.700 ;
        RECT 149.000 52.100 149.300 52.400 ;
        RECT 151.000 52.100 151.400 52.500 ;
        RECT 146.200 51.800 147.200 52.100 ;
        RECT 146.800 51.100 147.200 51.800 ;
        RECT 149.000 51.100 149.400 52.100 ;
        RECT 151.000 51.800 151.700 52.100 ;
        RECT 151.100 51.100 151.700 51.800 ;
        RECT 153.400 51.100 153.800 53.300 ;
        RECT 154.200 53.600 156.300 53.900 ;
        RECT 156.800 53.800 157.800 54.200 ;
        RECT 160.600 53.800 161.400 54.200 ;
        RECT 154.200 52.500 154.500 53.600 ;
        RECT 156.800 53.500 157.100 53.800 ;
        RECT 156.700 53.300 157.100 53.500 ;
        RECT 156.300 53.000 157.100 53.300 ;
        RECT 154.200 51.500 154.600 52.500 ;
        RECT 156.300 52.200 156.700 53.000 ;
        RECT 159.800 52.800 160.700 53.200 ;
        RECT 162.500 52.500 162.800 55.700 ;
        RECT 165.400 55.500 167.300 55.800 ;
        RECT 165.400 54.400 165.800 55.200 ;
        RECT 166.200 54.400 166.600 55.200 ;
        RECT 167.000 54.500 167.300 55.500 ;
        RECT 167.000 54.100 167.700 54.500 ;
        RECT 168.000 54.200 168.300 56.100 ;
        RECT 170.200 55.600 170.600 59.900 ;
        RECT 172.300 57.900 172.900 59.900 ;
        RECT 174.600 57.900 175.000 59.900 ;
        RECT 176.800 58.200 177.200 59.900 ;
        RECT 176.800 57.900 177.800 58.200 ;
        RECT 172.600 57.500 173.000 57.900 ;
        RECT 174.700 57.600 175.000 57.900 ;
        RECT 174.300 57.300 176.100 57.600 ;
        RECT 177.400 57.500 177.800 57.900 ;
        RECT 174.300 57.200 174.700 57.300 ;
        RECT 175.700 57.200 176.100 57.300 ;
        RECT 172.200 56.600 172.900 57.000 ;
        RECT 172.600 56.100 172.900 56.600 ;
        RECT 173.700 56.500 174.800 56.800 ;
        RECT 173.700 56.400 174.100 56.500 ;
        RECT 172.600 55.800 173.800 56.100 ;
        RECT 168.600 54.800 169.000 55.600 ;
        RECT 170.200 55.300 172.300 55.600 ;
        RECT 167.000 53.900 167.500 54.100 ;
        RECT 160.800 52.200 162.800 52.500 ;
        RECT 156.300 51.800 157.000 52.200 ;
        RECT 160.800 52.100 161.100 52.200 ;
        RECT 160.600 51.800 161.100 52.100 ;
        RECT 162.200 52.100 162.800 52.200 ;
        RECT 165.400 53.600 167.500 53.900 ;
        RECT 168.000 53.800 169.000 54.200 ;
        RECT 165.400 52.500 165.700 53.600 ;
        RECT 168.000 53.500 168.300 53.800 ;
        RECT 167.900 53.300 168.300 53.500 ;
        RECT 167.500 53.000 168.300 53.300 ;
        RECT 170.200 53.600 170.600 55.300 ;
        RECT 171.900 55.200 172.300 55.300 ;
        RECT 173.500 55.100 173.800 55.800 ;
        RECT 174.500 55.900 174.800 56.500 ;
        RECT 175.100 56.500 175.500 56.600 ;
        RECT 177.400 56.500 177.800 56.600 ;
        RECT 175.100 56.200 177.800 56.500 ;
        RECT 174.500 55.700 176.900 55.900 ;
        RECT 179.000 55.700 179.400 59.900 ;
        RECT 174.500 55.600 179.400 55.700 ;
        RECT 176.500 55.500 179.400 55.600 ;
        RECT 176.600 55.400 179.400 55.500 ;
        RECT 174.200 55.100 174.600 55.200 ;
        RECT 171.100 54.900 171.500 55.000 ;
        RECT 171.100 54.600 173.000 54.900 ;
        RECT 173.400 54.800 174.600 55.100 ;
        RECT 175.800 55.100 176.200 55.200 ;
        RECT 175.800 54.800 178.300 55.100 ;
        RECT 172.600 54.500 173.000 54.600 ;
        RECT 173.500 54.200 173.800 54.800 ;
        RECT 176.600 54.700 177.000 54.800 ;
        RECT 177.900 54.700 178.300 54.800 ;
        RECT 177.100 54.200 177.500 54.300 ;
        RECT 173.500 53.900 179.000 54.200 ;
        RECT 173.700 53.800 174.100 53.900 ;
        RECT 170.200 53.300 172.100 53.600 ;
        RECT 156.300 51.500 156.700 51.800 ;
        RECT 160.600 51.100 161.000 51.800 ;
        RECT 162.200 51.100 162.600 52.100 ;
        RECT 165.400 51.500 165.800 52.500 ;
        RECT 167.500 51.500 167.900 53.000 ;
        RECT 170.200 51.100 170.600 53.300 ;
        RECT 171.700 53.200 172.100 53.300 ;
        RECT 176.600 52.800 176.900 53.900 ;
        RECT 178.200 53.800 179.000 53.900 ;
        RECT 175.700 52.700 176.100 52.800 ;
        RECT 172.600 52.100 173.000 52.500 ;
        RECT 174.700 52.400 176.100 52.700 ;
        RECT 176.600 52.400 177.000 52.800 ;
        RECT 174.700 52.100 175.000 52.400 ;
        RECT 177.400 52.100 177.800 52.500 ;
        RECT 172.300 51.800 173.000 52.100 ;
        RECT 172.300 51.100 172.900 51.800 ;
        RECT 174.600 51.100 175.000 52.100 ;
        RECT 176.800 51.800 177.800 52.100 ;
        RECT 176.800 51.100 177.200 51.800 ;
        RECT 179.000 51.100 179.400 53.500 ;
        RECT 0.600 47.500 1.000 49.900 ;
        RECT 2.800 49.200 3.200 49.900 ;
        RECT 2.200 48.900 3.200 49.200 ;
        RECT 5.000 48.900 5.400 49.900 ;
        RECT 7.100 49.200 7.700 49.900 ;
        RECT 7.000 48.900 7.700 49.200 ;
        RECT 2.200 48.500 2.600 48.900 ;
        RECT 5.000 48.600 5.300 48.900 ;
        RECT 3.000 48.200 3.400 48.600 ;
        RECT 3.900 48.300 5.300 48.600 ;
        RECT 7.000 48.500 7.400 48.900 ;
        RECT 3.900 48.200 4.300 48.300 ;
        RECT 1.000 47.100 1.800 47.200 ;
        RECT 3.100 47.100 3.400 48.200 ;
        RECT 7.900 47.700 8.300 47.800 ;
        RECT 9.400 47.700 9.800 49.900 ;
        RECT 10.200 47.800 10.600 48.600 ;
        RECT 7.900 47.400 9.800 47.700 ;
        RECT 5.900 47.100 6.300 47.200 ;
        RECT 1.000 46.800 6.500 47.100 ;
        RECT 2.500 46.700 2.900 46.800 ;
        RECT 1.700 46.200 2.100 46.300 ;
        RECT 3.000 46.200 3.400 46.300 ;
        RECT 6.200 46.200 6.500 46.800 ;
        RECT 7.000 46.400 7.400 46.500 ;
        RECT 1.700 45.900 4.200 46.200 ;
        RECT 3.800 45.800 4.200 45.900 ;
        RECT 6.200 45.800 6.600 46.200 ;
        RECT 7.000 46.100 8.900 46.400 ;
        RECT 8.500 46.000 8.900 46.100 ;
        RECT 0.600 45.500 3.400 45.600 ;
        RECT 0.600 45.400 3.500 45.500 ;
        RECT 0.600 45.300 5.500 45.400 ;
        RECT 0.600 41.100 1.000 45.300 ;
        RECT 3.100 45.100 5.500 45.300 ;
        RECT 2.200 44.500 4.900 44.800 ;
        RECT 2.200 44.400 2.600 44.500 ;
        RECT 4.500 44.400 4.900 44.500 ;
        RECT 5.200 44.500 5.500 45.100 ;
        RECT 6.200 45.200 6.500 45.800 ;
        RECT 7.700 45.700 8.100 45.800 ;
        RECT 9.400 45.700 9.800 47.400 ;
        RECT 7.700 45.400 9.800 45.700 ;
        RECT 6.200 44.900 7.400 45.200 ;
        RECT 5.900 44.500 6.300 44.600 ;
        RECT 5.200 44.200 6.300 44.500 ;
        RECT 7.100 44.400 7.400 44.900 ;
        RECT 7.100 44.000 7.800 44.400 ;
        RECT 3.900 43.700 4.300 43.800 ;
        RECT 5.300 43.700 5.700 43.800 ;
        RECT 2.200 43.100 2.600 43.500 ;
        RECT 3.900 43.400 5.700 43.700 ;
        RECT 5.000 43.100 5.300 43.400 ;
        RECT 7.000 43.100 7.400 43.500 ;
        RECT 2.200 42.800 3.200 43.100 ;
        RECT 2.800 41.100 3.200 42.800 ;
        RECT 5.000 41.100 5.400 43.100 ;
        RECT 7.100 41.100 7.700 43.100 ;
        RECT 9.400 41.100 9.800 45.400 ;
        RECT 11.000 41.100 11.400 49.900 ;
        RECT 13.700 49.200 14.100 49.500 ;
        RECT 13.400 48.800 14.100 49.200 ;
        RECT 13.700 48.000 14.100 48.800 ;
        RECT 15.800 48.500 16.200 49.500 ;
        RECT 13.300 47.700 14.100 48.000 ;
        RECT 13.300 47.500 13.700 47.700 ;
        RECT 13.300 47.200 13.600 47.500 ;
        RECT 15.900 47.400 16.200 48.500 ;
        RECT 12.600 46.800 13.600 47.200 ;
        RECT 14.100 47.100 16.200 47.400 ;
        RECT 14.100 46.900 14.600 47.100 ;
        RECT 12.600 45.400 13.000 46.200 ;
        RECT 13.300 44.900 13.600 46.800 ;
        RECT 13.900 46.500 14.600 46.900 ;
        RECT 14.300 45.500 14.600 46.500 ;
        RECT 15.000 45.800 15.400 46.600 ;
        RECT 15.800 45.800 16.200 46.600 ;
        RECT 14.300 45.200 16.200 45.500 ;
        RECT 13.300 44.600 14.100 44.900 ;
        RECT 13.700 41.100 14.100 44.600 ;
        RECT 15.900 43.500 16.200 45.200 ;
        RECT 15.800 41.500 16.200 43.500 ;
        RECT 16.600 41.100 17.000 49.900 ;
        RECT 19.500 49.200 19.900 49.900 ;
        RECT 19.000 48.800 19.900 49.200 ;
        RECT 17.400 47.800 17.800 48.600 ;
        RECT 19.500 48.200 19.900 48.800 ;
        RECT 19.000 47.900 19.900 48.200 ;
        RECT 17.400 47.100 17.800 47.200 ;
        RECT 18.200 47.100 18.600 47.600 ;
        RECT 17.400 46.800 18.600 47.100 ;
        RECT 19.000 41.100 19.400 47.900 ;
        RECT 21.400 47.600 21.800 49.900 ;
        RECT 23.000 47.600 23.400 49.900 ;
        RECT 24.600 47.600 25.000 49.900 ;
        RECT 26.200 47.600 26.600 49.900 ;
        RECT 20.600 47.200 21.800 47.600 ;
        RECT 22.300 47.200 23.400 47.600 ;
        RECT 23.900 47.200 25.000 47.600 ;
        RECT 25.700 47.200 26.600 47.600 ;
        RECT 27.800 48.500 28.200 49.500 ;
        RECT 27.800 47.400 28.100 48.500 ;
        RECT 29.900 48.000 30.300 49.500 ;
        RECT 29.900 47.700 30.700 48.000 ;
        RECT 30.300 47.500 30.700 47.700 ;
        RECT 20.600 45.800 21.000 47.200 ;
        RECT 22.300 46.900 22.700 47.200 ;
        RECT 23.900 46.900 24.300 47.200 ;
        RECT 25.700 46.900 26.100 47.200 ;
        RECT 27.800 47.100 29.900 47.400 ;
        RECT 21.400 46.500 22.700 46.900 ;
        RECT 23.100 46.500 24.300 46.900 ;
        RECT 24.800 46.500 26.100 46.900 ;
        RECT 29.400 46.900 29.900 47.100 ;
        RECT 30.400 47.200 30.700 47.500 ;
        RECT 30.400 47.100 31.400 47.200 ;
        RECT 31.800 47.100 32.200 47.200 ;
        RECT 22.300 45.800 22.700 46.500 ;
        RECT 23.900 45.800 24.300 46.500 ;
        RECT 25.700 45.800 26.100 46.500 ;
        RECT 27.800 45.800 28.200 46.600 ;
        RECT 28.600 45.800 29.000 46.600 ;
        RECT 29.400 46.500 30.100 46.900 ;
        RECT 30.400 46.800 32.200 47.100 ;
        RECT 20.600 45.400 21.800 45.800 ;
        RECT 22.300 45.400 23.400 45.800 ;
        RECT 23.900 45.400 25.000 45.800 ;
        RECT 25.700 45.400 26.600 45.800 ;
        RECT 29.400 45.500 29.700 46.500 ;
        RECT 19.800 44.400 20.200 45.200 ;
        RECT 21.400 41.100 21.800 45.400 ;
        RECT 23.000 41.100 23.400 45.400 ;
        RECT 24.600 41.100 25.000 45.400 ;
        RECT 26.200 41.100 26.600 45.400 ;
        RECT 27.800 45.200 29.700 45.500 ;
        RECT 27.800 43.500 28.100 45.200 ;
        RECT 30.400 44.900 30.700 46.800 ;
        RECT 31.000 46.100 31.400 46.200 ;
        RECT 32.600 46.100 33.000 49.900 ;
        RECT 33.400 48.100 33.800 48.600 ;
        RECT 35.000 48.100 35.400 48.200 ;
        RECT 33.400 47.800 35.400 48.100 ;
        RECT 35.800 47.500 36.200 49.900 ;
        RECT 38.000 49.200 38.400 49.900 ;
        RECT 37.400 48.900 38.400 49.200 ;
        RECT 40.200 48.900 40.600 49.900 ;
        RECT 42.300 49.200 42.900 49.900 ;
        RECT 42.200 48.900 42.900 49.200 ;
        RECT 37.400 48.500 37.800 48.900 ;
        RECT 40.200 48.600 40.500 48.900 ;
        RECT 38.200 48.200 38.600 48.600 ;
        RECT 39.100 48.300 40.500 48.600 ;
        RECT 42.200 48.500 42.600 48.900 ;
        RECT 39.100 48.200 39.500 48.300 ;
        RECT 36.200 47.100 37.000 47.200 ;
        RECT 38.300 47.100 38.600 48.200 ;
        RECT 43.100 47.700 43.500 47.800 ;
        RECT 44.600 47.700 45.000 49.900 ;
        RECT 43.100 47.400 45.000 47.700 ;
        RECT 41.100 47.100 41.500 47.200 ;
        RECT 36.200 46.800 41.700 47.100 ;
        RECT 37.700 46.700 38.100 46.800 ;
        RECT 31.000 45.800 33.000 46.100 ;
        RECT 36.900 46.200 37.300 46.300 ;
        RECT 38.200 46.200 38.600 46.300 ;
        RECT 36.900 45.900 39.400 46.200 ;
        RECT 39.000 45.800 39.400 45.900 ;
        RECT 31.000 45.400 31.400 45.800 ;
        RECT 29.900 44.600 30.700 44.900 ;
        RECT 27.800 41.500 28.200 43.500 ;
        RECT 29.900 41.100 30.300 44.600 ;
        RECT 32.600 41.100 33.000 45.800 ;
        RECT 35.800 45.500 38.600 45.600 ;
        RECT 35.800 45.400 38.700 45.500 ;
        RECT 35.800 45.300 40.700 45.400 ;
        RECT 35.800 41.100 36.200 45.300 ;
        RECT 38.300 45.100 40.700 45.300 ;
        RECT 37.400 44.500 40.100 44.800 ;
        RECT 37.400 44.400 37.800 44.500 ;
        RECT 39.700 44.400 40.100 44.500 ;
        RECT 40.400 44.500 40.700 45.100 ;
        RECT 41.400 45.200 41.700 46.800 ;
        RECT 42.200 46.400 42.600 46.500 ;
        RECT 42.200 46.100 44.100 46.400 ;
        RECT 43.700 46.000 44.100 46.100 ;
        RECT 42.900 45.700 43.300 45.800 ;
        RECT 44.600 45.700 45.000 47.400 ;
        RECT 46.200 47.600 46.600 49.900 ;
        RECT 47.800 47.600 48.200 49.900 ;
        RECT 49.400 47.600 49.800 49.900 ;
        RECT 51.000 47.600 51.400 49.900 ;
        RECT 53.400 48.800 53.800 49.900 ;
        RECT 52.600 47.800 53.000 48.600 ;
        RECT 46.200 47.200 47.100 47.600 ;
        RECT 47.800 47.200 48.900 47.600 ;
        RECT 49.400 47.200 50.500 47.600 ;
        RECT 51.000 47.200 52.200 47.600 ;
        RECT 53.500 47.200 53.800 48.800 ;
        RECT 55.100 48.200 55.500 48.600 ;
        RECT 55.000 47.800 55.400 48.200 ;
        RECT 55.800 47.900 56.200 49.900 ;
        RECT 46.700 46.900 47.100 47.200 ;
        RECT 48.500 46.900 48.900 47.200 ;
        RECT 50.100 46.900 50.500 47.200 ;
        RECT 46.700 46.500 48.000 46.900 ;
        RECT 48.500 46.500 49.700 46.900 ;
        RECT 50.100 46.500 51.400 46.900 ;
        RECT 46.700 45.800 47.100 46.500 ;
        RECT 48.500 45.800 48.900 46.500 ;
        RECT 50.100 45.800 50.500 46.500 ;
        RECT 51.800 45.800 52.200 47.200 ;
        RECT 53.400 46.800 53.800 47.200 ;
        RECT 42.900 45.400 45.000 45.700 ;
        RECT 41.400 44.900 42.600 45.200 ;
        RECT 41.100 44.500 41.500 44.600 ;
        RECT 40.400 44.200 41.500 44.500 ;
        RECT 42.300 44.400 42.600 44.900 ;
        RECT 42.300 44.000 43.000 44.400 ;
        RECT 39.100 43.700 39.500 43.800 ;
        RECT 40.500 43.700 40.900 43.800 ;
        RECT 37.400 43.100 37.800 43.500 ;
        RECT 39.100 43.400 40.900 43.700 ;
        RECT 40.200 43.100 40.500 43.400 ;
        RECT 42.200 43.100 42.600 43.500 ;
        RECT 37.400 42.800 38.400 43.100 ;
        RECT 38.000 41.100 38.400 42.800 ;
        RECT 40.200 41.100 40.600 43.100 ;
        RECT 42.300 41.100 42.900 43.100 ;
        RECT 44.600 41.100 45.000 45.400 ;
        RECT 46.200 45.400 47.100 45.800 ;
        RECT 47.800 45.400 48.900 45.800 ;
        RECT 49.400 45.400 50.500 45.800 ;
        RECT 51.000 45.400 52.200 45.800 ;
        RECT 46.200 41.100 46.600 45.400 ;
        RECT 47.800 41.100 48.200 45.400 ;
        RECT 49.400 41.100 49.800 45.400 ;
        RECT 51.000 41.100 51.400 45.400 ;
        RECT 53.500 45.100 53.800 46.800 ;
        RECT 54.200 45.400 54.600 46.200 ;
        RECT 55.000 46.100 55.400 46.200 ;
        RECT 55.900 46.100 56.200 47.900 ;
        RECT 59.000 48.900 59.400 49.900 ;
        RECT 63.000 48.900 63.400 49.900 ;
        RECT 64.600 49.200 65.000 49.900 ;
        RECT 59.000 47.200 59.300 48.900 ;
        RECT 62.800 48.800 63.400 48.900 ;
        RECT 64.500 48.800 65.000 49.200 ;
        RECT 68.300 49.200 68.700 49.900 ;
        RECT 68.300 48.800 69.000 49.200 ;
        RECT 59.800 47.800 60.200 48.600 ;
        RECT 62.800 48.500 64.800 48.800 ;
        RECT 56.600 47.100 57.000 47.200 ;
        RECT 58.200 47.100 58.600 47.200 ;
        RECT 56.600 46.800 58.600 47.100 ;
        RECT 59.000 47.100 59.400 47.200 ;
        RECT 60.600 47.100 61.000 47.200 ;
        RECT 59.000 46.800 61.000 47.100 ;
        RECT 56.600 46.400 57.000 46.800 ;
        RECT 57.400 46.100 57.800 46.200 ;
        RECT 55.000 45.800 56.200 46.100 ;
        RECT 57.000 45.800 57.800 46.100 ;
        RECT 55.100 45.100 55.400 45.800 ;
        RECT 57.000 45.600 57.400 45.800 ;
        RECT 58.200 45.400 58.600 46.200 ;
        RECT 59.000 45.100 59.300 46.800 ;
        RECT 62.800 45.200 63.100 48.500 ;
        RECT 68.300 48.200 68.700 48.800 ;
        RECT 67.800 47.900 68.700 48.200 ;
        RECT 64.200 46.800 65.000 47.200 ;
        RECT 63.400 46.100 64.200 46.200 ;
        RECT 66.200 46.100 66.600 46.200 ;
        RECT 63.400 45.800 66.600 46.100 ;
        RECT 53.400 44.700 54.300 45.100 ;
        RECT 53.900 41.100 54.300 44.700 ;
        RECT 55.000 41.100 55.400 45.100 ;
        RECT 55.800 44.800 57.800 45.100 ;
        RECT 55.800 41.100 56.200 44.800 ;
        RECT 57.400 41.100 57.800 44.800 ;
        RECT 58.500 44.700 59.400 45.100 ;
        RECT 61.400 44.900 63.100 45.200 ;
        RECT 61.400 44.800 61.800 44.900 ;
        RECT 58.500 41.100 58.900 44.700 ;
        RECT 61.500 44.500 61.800 44.800 ;
        RECT 62.300 44.500 64.100 44.600 ;
        RECT 60.600 41.500 61.000 44.500 ;
        RECT 61.400 41.700 61.800 44.500 ;
        RECT 62.200 44.300 64.100 44.500 ;
        RECT 60.700 41.400 61.000 41.500 ;
        RECT 62.200 41.500 62.600 44.300 ;
        RECT 63.800 44.100 64.100 44.300 ;
        RECT 64.700 44.400 66.500 44.700 ;
        RECT 64.700 44.100 65.000 44.400 ;
        RECT 62.200 41.400 62.500 41.500 ;
        RECT 60.700 41.100 62.500 41.400 ;
        RECT 63.000 41.400 63.400 44.000 ;
        RECT 63.800 41.700 64.200 44.100 ;
        RECT 64.600 41.400 65.000 44.100 ;
        RECT 63.000 41.100 65.000 41.400 ;
        RECT 66.200 44.100 66.500 44.400 ;
        RECT 66.200 41.100 66.600 44.100 ;
        RECT 67.800 41.100 68.200 47.900 ;
        RECT 69.400 47.100 69.800 49.900 ;
        RECT 71.000 47.500 71.400 49.900 ;
        RECT 73.200 49.200 73.600 49.900 ;
        RECT 72.600 48.900 73.600 49.200 ;
        RECT 75.400 48.900 75.800 49.900 ;
        RECT 77.500 49.200 78.100 49.900 ;
        RECT 77.400 48.900 78.100 49.200 ;
        RECT 72.600 48.500 73.000 48.900 ;
        RECT 75.400 48.600 75.700 48.900 ;
        RECT 73.400 48.200 73.800 48.600 ;
        RECT 74.300 48.300 75.700 48.600 ;
        RECT 77.400 48.500 77.800 48.900 ;
        RECT 74.300 48.200 74.700 48.300 ;
        RECT 68.600 46.800 69.800 47.100 ;
        RECT 71.400 47.100 72.200 47.200 ;
        RECT 73.500 47.100 73.800 48.200 ;
        RECT 76.600 47.800 77.000 48.200 ;
        RECT 76.600 47.200 76.900 47.800 ;
        RECT 78.300 47.700 78.700 47.800 ;
        RECT 79.800 47.700 80.200 49.900 ;
        RECT 78.300 47.400 80.200 47.700 ;
        RECT 80.600 47.500 81.000 49.900 ;
        RECT 82.800 49.200 83.200 49.900 ;
        RECT 82.200 48.900 83.200 49.200 ;
        RECT 85.000 48.900 85.400 49.900 ;
        RECT 87.100 49.200 87.700 49.900 ;
        RECT 87.000 48.900 87.700 49.200 ;
        RECT 89.400 49.100 89.800 49.900 ;
        RECT 90.200 49.100 90.600 49.200 ;
        RECT 82.200 48.500 82.600 48.900 ;
        RECT 85.000 48.600 85.300 48.900 ;
        RECT 83.000 48.200 83.400 48.600 ;
        RECT 83.900 48.300 85.300 48.600 ;
        RECT 87.000 48.500 87.400 48.900 ;
        RECT 89.400 48.800 90.600 49.100 ;
        RECT 83.900 48.200 84.300 48.300 ;
        RECT 76.300 47.100 76.900 47.200 ;
        RECT 71.400 46.800 76.900 47.100 ;
        RECT 68.600 46.200 68.900 46.800 ;
        RECT 68.600 45.800 69.000 46.200 ;
        RECT 68.600 45.100 69.000 45.200 ;
        RECT 69.400 45.100 69.800 46.800 ;
        RECT 72.900 46.700 73.300 46.800 ;
        RECT 72.100 46.200 72.500 46.300 ;
        RECT 72.100 46.100 74.600 46.200 ;
        RECT 75.000 46.100 75.400 46.200 ;
        RECT 72.100 45.900 75.400 46.100 ;
        RECT 74.200 45.800 75.400 45.900 ;
        RECT 68.600 44.800 69.800 45.100 ;
        RECT 68.600 44.400 69.000 44.800 ;
        RECT 69.400 41.100 69.800 44.800 ;
        RECT 71.000 45.500 73.800 45.600 ;
        RECT 71.000 45.400 73.900 45.500 ;
        RECT 71.000 45.300 75.900 45.400 ;
        RECT 71.000 41.100 71.400 45.300 ;
        RECT 73.500 45.100 75.900 45.300 ;
        RECT 72.600 44.500 75.300 44.800 ;
        RECT 72.600 44.400 73.000 44.500 ;
        RECT 74.900 44.400 75.300 44.500 ;
        RECT 75.600 44.500 75.900 45.100 ;
        RECT 76.600 45.200 76.900 46.800 ;
        RECT 77.400 46.400 77.800 46.500 ;
        RECT 77.400 46.100 79.300 46.400 ;
        RECT 78.900 46.000 79.300 46.100 ;
        RECT 78.100 45.700 78.500 45.800 ;
        RECT 79.800 45.700 80.200 47.400 ;
        RECT 81.000 47.100 81.800 47.200 ;
        RECT 83.100 47.100 83.400 48.200 ;
        RECT 87.900 47.700 88.300 47.800 ;
        RECT 89.400 47.700 89.800 48.800 ;
        RECT 87.900 47.400 89.800 47.700 ;
        RECT 85.900 47.100 86.300 47.200 ;
        RECT 81.000 46.800 86.500 47.100 ;
        RECT 82.500 46.700 82.900 46.800 ;
        RECT 81.700 46.200 82.100 46.300 ;
        RECT 81.700 45.900 84.200 46.200 ;
        RECT 83.800 45.800 84.200 45.900 ;
        RECT 78.100 45.400 80.200 45.700 ;
        RECT 76.600 44.900 77.800 45.200 ;
        RECT 76.300 44.500 76.700 44.600 ;
        RECT 75.600 44.200 76.700 44.500 ;
        RECT 77.500 44.400 77.800 44.900 ;
        RECT 77.500 44.000 78.200 44.400 ;
        RECT 74.300 43.700 74.700 43.800 ;
        RECT 75.700 43.700 76.100 43.800 ;
        RECT 72.600 43.100 73.000 43.500 ;
        RECT 74.300 43.400 76.100 43.700 ;
        RECT 75.400 43.100 75.700 43.400 ;
        RECT 77.400 43.100 77.800 43.500 ;
        RECT 72.600 42.800 73.600 43.100 ;
        RECT 73.200 41.100 73.600 42.800 ;
        RECT 75.400 41.100 75.800 43.100 ;
        RECT 77.500 41.100 78.100 43.100 ;
        RECT 79.800 41.100 80.200 45.400 ;
        RECT 80.600 45.500 83.400 45.600 ;
        RECT 80.600 45.400 83.500 45.500 ;
        RECT 80.600 45.300 85.500 45.400 ;
        RECT 80.600 41.100 81.000 45.300 ;
        RECT 83.100 45.100 85.500 45.300 ;
        RECT 82.200 44.500 84.900 44.800 ;
        RECT 82.200 44.400 82.600 44.500 ;
        RECT 84.500 44.400 84.900 44.500 ;
        RECT 85.200 44.500 85.500 45.100 ;
        RECT 86.200 45.200 86.500 46.800 ;
        RECT 87.000 46.400 87.400 46.500 ;
        RECT 87.000 46.100 88.900 46.400 ;
        RECT 88.500 46.000 88.900 46.100 ;
        RECT 87.700 45.700 88.100 45.800 ;
        RECT 89.400 45.700 89.800 47.400 ;
        RECT 91.800 48.500 92.200 49.500 ;
        RECT 91.800 47.400 92.100 48.500 ;
        RECT 93.900 48.200 94.300 49.500 ;
        RECT 93.400 48.000 94.300 48.200 ;
        RECT 93.400 47.800 94.700 48.000 ;
        RECT 93.900 47.700 94.700 47.800 ;
        RECT 94.300 47.500 94.700 47.700 ;
        RECT 91.800 47.100 93.900 47.400 ;
        RECT 93.400 46.900 93.900 47.100 ;
        RECT 94.400 47.200 94.700 47.500 ;
        RECT 91.800 45.800 92.200 46.600 ;
        RECT 92.600 45.800 93.000 46.600 ;
        RECT 93.400 46.500 94.100 46.900 ;
        RECT 94.400 46.800 95.400 47.200 ;
        RECT 87.700 45.400 89.800 45.700 ;
        RECT 93.400 45.500 93.700 46.500 ;
        RECT 86.200 44.900 87.400 45.200 ;
        RECT 85.900 44.500 86.300 44.600 ;
        RECT 85.200 44.200 86.300 44.500 ;
        RECT 87.100 44.400 87.400 44.900 ;
        RECT 87.100 44.200 87.800 44.400 ;
        RECT 87.100 44.000 88.200 44.200 ;
        RECT 87.500 43.800 88.200 44.000 ;
        RECT 83.900 43.700 84.300 43.800 ;
        RECT 85.300 43.700 85.700 43.800 ;
        RECT 82.200 43.100 82.600 43.500 ;
        RECT 83.900 43.400 85.700 43.700 ;
        RECT 85.000 43.100 85.300 43.400 ;
        RECT 87.000 43.100 87.400 43.500 ;
        RECT 82.200 42.800 83.200 43.100 ;
        RECT 82.800 41.100 83.200 42.800 ;
        RECT 85.000 41.100 85.400 43.100 ;
        RECT 87.100 41.100 87.700 43.100 ;
        RECT 89.400 41.100 89.800 45.400 ;
        RECT 91.800 45.200 93.700 45.500 ;
        RECT 91.800 43.500 92.100 45.200 ;
        RECT 94.400 44.900 94.700 46.800 ;
        RECT 95.000 46.100 95.400 46.200 ;
        RECT 96.600 46.100 97.000 49.900 ;
        RECT 99.700 49.200 100.500 49.900 ;
        RECT 99.700 48.800 101.000 49.200 ;
        RECT 97.400 47.800 97.800 48.600 ;
        RECT 99.700 47.900 100.500 48.800 ;
        RECT 103.700 47.900 104.500 49.900 ;
        RECT 99.000 46.400 99.400 47.200 ;
        RECT 99.900 46.200 100.200 47.900 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 101.400 47.100 101.800 47.200 ;
        RECT 103.000 47.100 103.400 47.200 ;
        RECT 101.400 46.800 103.400 47.100 ;
        RECT 100.600 46.600 100.900 46.800 ;
        RECT 100.500 46.200 100.900 46.600 ;
        RECT 103.000 46.400 103.400 46.800 ;
        RECT 103.900 46.200 104.200 47.900 ;
        RECT 104.600 46.800 105.000 47.200 ;
        RECT 106.200 46.800 106.600 47.600 ;
        RECT 104.600 46.600 104.900 46.800 ;
        RECT 104.500 46.200 104.900 46.600 ;
        RECT 95.000 45.800 97.000 46.100 ;
        RECT 98.200 46.100 98.600 46.200 ;
        RECT 98.200 45.800 99.000 46.100 ;
        RECT 99.800 45.800 100.200 46.200 ;
        RECT 95.000 45.400 95.400 45.800 ;
        RECT 93.900 44.600 94.700 44.900 ;
        RECT 91.800 41.500 92.200 43.500 ;
        RECT 93.900 41.100 94.300 44.600 ;
        RECT 96.600 41.100 97.000 45.800 ;
        RECT 98.600 45.600 99.000 45.800 ;
        RECT 99.900 45.700 100.200 45.800 ;
        RECT 99.900 45.400 100.900 45.700 ;
        RECT 101.400 45.400 101.800 46.200 ;
        RECT 102.200 46.100 102.600 46.200 ;
        RECT 102.200 45.800 103.000 46.100 ;
        RECT 103.800 45.800 104.200 46.200 ;
        RECT 102.600 45.600 103.000 45.800 ;
        RECT 103.900 45.700 104.200 45.800 ;
        RECT 103.900 45.400 104.900 45.700 ;
        RECT 105.400 45.400 105.800 46.200 ;
        RECT 100.600 45.100 100.900 45.400 ;
        RECT 104.600 45.100 104.900 45.400 ;
        RECT 98.200 44.800 100.200 45.100 ;
        RECT 98.200 41.100 98.600 44.800 ;
        RECT 99.800 41.400 100.200 44.800 ;
        RECT 100.600 41.700 101.000 45.100 ;
        RECT 101.400 41.400 101.800 45.100 ;
        RECT 99.800 41.100 101.800 41.400 ;
        RECT 102.200 44.800 104.200 45.100 ;
        RECT 102.200 41.100 102.600 44.800 ;
        RECT 103.800 41.400 104.200 44.800 ;
        RECT 104.600 41.700 105.000 45.100 ;
        RECT 105.400 41.400 105.800 45.100 ;
        RECT 103.800 41.100 105.800 41.400 ;
        RECT 107.000 41.100 107.400 49.900 ;
        RECT 107.800 47.800 108.200 48.600 ;
        RECT 108.600 41.100 109.000 49.900 ;
        RECT 109.400 47.500 109.800 49.900 ;
        RECT 111.600 49.200 112.000 49.900 ;
        RECT 111.000 48.900 112.000 49.200 ;
        RECT 113.800 48.900 114.200 49.900 ;
        RECT 115.900 49.200 116.500 49.900 ;
        RECT 115.800 48.900 116.500 49.200 ;
        RECT 111.000 48.500 111.400 48.900 ;
        RECT 113.800 48.600 114.100 48.900 ;
        RECT 111.800 48.200 112.200 48.600 ;
        RECT 112.700 48.300 114.100 48.600 ;
        RECT 115.800 48.500 116.200 48.900 ;
        RECT 112.700 48.200 113.100 48.300 ;
        RECT 109.800 47.100 110.600 47.200 ;
        RECT 111.900 47.100 112.200 48.200 ;
        RECT 116.700 47.700 117.100 47.800 ;
        RECT 118.200 47.700 118.600 49.900 ;
        RECT 119.000 47.900 119.400 49.900 ;
        RECT 119.800 48.000 120.200 49.900 ;
        RECT 121.400 48.000 121.800 49.900 ;
        RECT 119.800 47.900 121.800 48.000 ;
        RECT 116.700 47.400 118.600 47.700 ;
        RECT 114.700 47.100 115.100 47.200 ;
        RECT 109.800 46.800 115.300 47.100 ;
        RECT 111.300 46.700 111.700 46.800 ;
        RECT 110.500 46.200 110.900 46.300 ;
        RECT 110.500 45.900 113.000 46.200 ;
        RECT 112.600 45.800 113.000 45.900 ;
        RECT 109.400 45.500 112.200 45.600 ;
        RECT 109.400 45.400 112.300 45.500 ;
        RECT 109.400 45.300 114.300 45.400 ;
        RECT 109.400 41.100 109.800 45.300 ;
        RECT 111.900 45.100 114.300 45.300 ;
        RECT 111.000 44.500 113.700 44.800 ;
        RECT 111.000 44.400 111.400 44.500 ;
        RECT 113.300 44.400 113.700 44.500 ;
        RECT 114.000 44.500 114.300 45.100 ;
        RECT 115.000 45.200 115.300 46.800 ;
        RECT 115.800 46.400 116.200 46.500 ;
        RECT 115.800 46.100 117.700 46.400 ;
        RECT 117.300 46.000 117.700 46.100 ;
        RECT 116.500 45.700 116.900 45.800 ;
        RECT 118.200 45.700 118.600 47.400 ;
        RECT 119.100 47.200 119.400 47.900 ;
        RECT 119.900 47.700 121.700 47.900 ;
        RECT 122.200 47.800 122.600 48.600 ;
        RECT 121.000 47.200 121.400 47.400 ;
        RECT 119.000 46.800 120.300 47.200 ;
        RECT 121.000 46.900 121.800 47.200 ;
        RECT 121.400 46.800 121.800 46.900 ;
        RECT 116.500 45.400 118.600 45.700 ;
        RECT 115.000 44.900 116.200 45.200 ;
        RECT 114.700 44.500 115.100 44.600 ;
        RECT 114.000 44.200 115.100 44.500 ;
        RECT 115.900 44.400 116.200 44.900 ;
        RECT 115.900 44.000 116.600 44.400 ;
        RECT 112.700 43.700 113.100 43.800 ;
        RECT 114.100 43.700 114.500 43.800 ;
        RECT 111.000 43.100 111.400 43.500 ;
        RECT 112.700 43.400 114.500 43.700 ;
        RECT 113.800 43.100 114.100 43.400 ;
        RECT 115.800 43.100 116.200 43.500 ;
        RECT 111.000 42.800 112.000 43.100 ;
        RECT 111.600 41.100 112.000 42.800 ;
        RECT 113.800 41.100 114.200 43.100 ;
        RECT 115.900 41.100 116.500 43.100 ;
        RECT 118.200 41.100 118.600 45.400 ;
        RECT 119.000 45.100 119.400 45.200 ;
        RECT 120.000 45.100 120.300 46.800 ;
        RECT 120.600 45.800 121.000 46.600 ;
        RECT 123.000 46.100 123.400 49.900 ;
        RECT 123.800 48.000 124.200 49.900 ;
        RECT 125.400 48.000 125.800 49.900 ;
        RECT 123.800 47.900 125.800 48.000 ;
        RECT 126.200 47.900 126.600 49.900 ;
        RECT 128.900 48.000 129.300 49.500 ;
        RECT 131.000 48.500 131.400 49.500 ;
        RECT 123.900 47.700 125.700 47.900 ;
        RECT 124.200 47.200 124.600 47.400 ;
        RECT 126.200 47.200 126.500 47.900 ;
        RECT 128.500 47.700 129.300 48.000 ;
        RECT 128.500 47.500 128.900 47.700 ;
        RECT 128.500 47.200 128.800 47.500 ;
        RECT 131.100 47.400 131.400 48.500 ;
        RECT 131.800 47.800 132.200 48.600 ;
        RECT 123.800 46.900 124.600 47.200 ;
        RECT 123.800 46.800 124.200 46.900 ;
        RECT 125.300 46.800 126.600 47.200 ;
        RECT 127.000 47.100 127.400 47.200 ;
        RECT 127.800 47.100 128.800 47.200 ;
        RECT 127.000 46.800 128.800 47.100 ;
        RECT 129.300 47.100 131.400 47.400 ;
        RECT 129.300 46.900 129.800 47.100 ;
        RECT 124.600 46.100 125.000 46.600 ;
        RECT 123.000 45.800 125.000 46.100 ;
        RECT 119.000 44.800 119.700 45.100 ;
        RECT 120.000 44.800 120.500 45.100 ;
        RECT 119.400 44.200 119.700 44.800 ;
        RECT 119.400 43.800 119.800 44.200 ;
        RECT 120.100 41.100 120.500 44.800 ;
        RECT 123.000 41.100 123.400 45.800 ;
        RECT 125.300 45.100 125.600 46.800 ;
        RECT 127.800 45.400 128.200 46.200 ;
        RECT 126.200 45.100 126.600 45.200 ;
        RECT 125.100 44.800 125.600 45.100 ;
        RECT 125.900 44.800 126.600 45.100 ;
        RECT 128.500 44.900 128.800 46.800 ;
        RECT 129.100 46.500 129.800 46.900 ;
        RECT 129.500 45.500 129.800 46.500 ;
        RECT 130.200 45.800 130.600 46.600 ;
        RECT 131.000 45.800 131.400 46.600 ;
        RECT 129.500 45.200 131.400 45.500 ;
        RECT 125.100 41.100 125.500 44.800 ;
        RECT 125.900 44.200 126.200 44.800 ;
        RECT 128.500 44.600 129.300 44.900 ;
        RECT 125.800 43.800 126.200 44.200 ;
        RECT 128.900 41.100 129.300 44.600 ;
        RECT 131.100 43.500 131.400 45.200 ;
        RECT 131.000 41.500 131.400 43.500 ;
        RECT 132.600 41.100 133.000 49.900 ;
        RECT 133.400 48.500 133.800 49.500 ;
        RECT 133.400 47.400 133.700 48.500 ;
        RECT 135.500 48.000 135.900 49.500 ;
        RECT 135.500 47.700 136.300 48.000 ;
        RECT 135.900 47.500 136.300 47.700 ;
        RECT 133.400 47.100 135.500 47.400 ;
        RECT 135.000 46.900 135.500 47.100 ;
        RECT 136.000 47.200 136.300 47.500 ;
        RECT 133.400 45.800 133.800 46.600 ;
        RECT 134.200 45.800 134.600 46.600 ;
        RECT 135.000 46.500 135.700 46.900 ;
        RECT 136.000 46.800 137.000 47.200 ;
        RECT 135.000 45.500 135.300 46.500 ;
        RECT 133.400 45.200 135.300 45.500 ;
        RECT 133.400 43.500 133.700 45.200 ;
        RECT 136.000 44.900 136.300 46.800 ;
        RECT 136.600 46.100 137.000 46.200 ;
        RECT 138.200 46.100 138.600 49.900 ;
        RECT 139.000 48.100 139.400 48.600 ;
        RECT 140.600 48.100 141.000 48.200 ;
        RECT 139.000 47.800 141.000 48.100 ;
        RECT 142.200 47.600 142.600 49.900 ;
        RECT 143.800 47.600 144.200 49.900 ;
        RECT 145.400 47.600 145.800 49.900 ;
        RECT 147.000 47.600 147.400 49.900 ;
        RECT 136.600 45.800 138.600 46.100 ;
        RECT 136.600 45.400 137.000 45.800 ;
        RECT 135.500 44.600 136.300 44.900 ;
        RECT 133.400 41.500 133.800 43.500 ;
        RECT 135.500 42.200 135.900 44.600 ;
        RECT 135.500 41.800 136.200 42.200 ;
        RECT 135.500 41.100 135.900 41.800 ;
        RECT 138.200 41.100 138.600 45.800 ;
        RECT 141.400 47.200 142.600 47.600 ;
        RECT 143.100 47.200 144.200 47.600 ;
        RECT 144.700 47.200 145.800 47.600 ;
        RECT 146.500 47.200 147.400 47.600 ;
        RECT 148.600 48.500 149.000 49.500 ;
        RECT 148.600 47.400 148.900 48.500 ;
        RECT 150.700 48.000 151.100 49.500 ;
        RECT 153.400 48.000 153.800 49.900 ;
        RECT 155.000 48.000 155.400 49.900 ;
        RECT 150.700 47.700 151.500 48.000 ;
        RECT 153.400 47.900 155.400 48.000 ;
        RECT 155.800 47.900 156.200 49.900 ;
        RECT 153.500 47.700 155.300 47.900 ;
        RECT 151.100 47.500 151.500 47.700 ;
        RECT 141.400 45.800 141.800 47.200 ;
        RECT 143.100 46.900 143.500 47.200 ;
        RECT 144.700 46.900 145.100 47.200 ;
        RECT 146.500 46.900 146.900 47.200 ;
        RECT 148.600 47.100 150.700 47.400 ;
        RECT 142.200 46.500 143.500 46.900 ;
        RECT 143.900 46.500 145.100 46.900 ;
        RECT 145.600 46.500 146.900 46.900 ;
        RECT 150.200 46.900 150.700 47.100 ;
        RECT 151.200 47.200 151.500 47.500 ;
        RECT 153.800 47.200 154.200 47.400 ;
        RECT 155.800 47.200 156.100 47.900 ;
        RECT 156.600 47.700 157.000 49.900 ;
        RECT 158.700 49.200 159.300 49.900 ;
        RECT 158.700 48.900 159.400 49.200 ;
        RECT 161.000 48.900 161.400 49.900 ;
        RECT 163.200 49.200 163.600 49.900 ;
        RECT 163.200 48.900 164.200 49.200 ;
        RECT 159.000 48.500 159.400 48.900 ;
        RECT 161.100 48.600 161.400 48.900 ;
        RECT 161.100 48.300 162.500 48.600 ;
        RECT 162.100 48.200 162.500 48.300 ;
        RECT 163.000 48.200 163.400 48.600 ;
        RECT 163.800 48.500 164.200 48.900 ;
        RECT 158.100 47.700 158.500 47.800 ;
        RECT 156.600 47.400 158.500 47.700 ;
        RECT 143.100 45.800 143.500 46.500 ;
        RECT 144.700 45.800 145.100 46.500 ;
        RECT 146.500 45.800 146.900 46.500 ;
        RECT 148.600 45.800 149.000 46.600 ;
        RECT 149.400 45.800 149.800 46.600 ;
        RECT 150.200 46.500 150.900 46.900 ;
        RECT 151.200 46.800 152.200 47.200 ;
        RECT 153.400 46.900 154.200 47.200 ;
        RECT 153.400 46.800 153.800 46.900 ;
        RECT 154.900 46.800 156.200 47.200 ;
        RECT 141.400 45.400 142.600 45.800 ;
        RECT 143.100 45.400 144.200 45.800 ;
        RECT 144.700 45.400 145.800 45.800 ;
        RECT 146.500 45.400 147.400 45.800 ;
        RECT 150.200 45.500 150.500 46.500 ;
        RECT 142.200 41.100 142.600 45.400 ;
        RECT 143.800 41.100 144.200 45.400 ;
        RECT 145.400 41.100 145.800 45.400 ;
        RECT 147.000 41.100 147.400 45.400 ;
        RECT 148.600 45.200 150.500 45.500 ;
        RECT 148.600 43.500 148.900 45.200 ;
        RECT 151.200 44.900 151.500 46.800 ;
        RECT 151.800 45.400 152.200 46.200 ;
        RECT 154.200 45.800 154.600 46.600 ;
        RECT 154.900 45.100 155.200 46.800 ;
        RECT 156.600 45.700 157.000 47.400 ;
        RECT 160.100 47.100 160.500 47.200 ;
        RECT 163.000 47.100 163.300 48.200 ;
        RECT 165.400 47.500 165.800 49.900 ;
        RECT 166.200 48.000 166.600 49.900 ;
        RECT 167.800 48.000 168.200 49.900 ;
        RECT 166.200 47.900 168.200 48.000 ;
        RECT 168.600 47.900 169.000 49.900 ;
        RECT 166.300 47.700 168.100 47.900 ;
        RECT 166.600 47.200 167.000 47.400 ;
        RECT 168.600 47.200 168.900 47.900 ;
        RECT 164.600 47.100 165.400 47.200 ;
        RECT 159.900 46.800 165.400 47.100 ;
        RECT 166.200 46.900 167.000 47.200 ;
        RECT 166.200 46.800 166.600 46.900 ;
        RECT 167.700 46.800 169.000 47.200 ;
        RECT 159.000 46.400 159.400 46.500 ;
        RECT 157.500 46.100 159.400 46.400 ;
        RECT 159.900 46.200 160.200 46.800 ;
        RECT 163.500 46.700 163.900 46.800 ;
        RECT 164.300 46.200 164.700 46.300 ;
        RECT 157.500 46.000 157.900 46.100 ;
        RECT 159.800 45.800 160.200 46.200 ;
        RECT 161.400 46.100 161.800 46.200 ;
        RECT 162.200 46.100 164.700 46.200 ;
        RECT 161.400 45.900 164.700 46.100 ;
        RECT 161.400 45.800 162.600 45.900 ;
        RECT 167.000 45.800 167.400 46.600 ;
        RECT 158.300 45.700 158.700 45.800 ;
        RECT 156.600 45.400 158.700 45.700 ;
        RECT 155.800 45.100 156.200 45.200 ;
        RECT 150.700 44.600 151.500 44.900 ;
        RECT 154.700 44.800 155.200 45.100 ;
        RECT 155.500 44.800 156.200 45.100 ;
        RECT 148.600 41.500 149.000 43.500 ;
        RECT 150.700 42.200 151.100 44.600 ;
        RECT 150.700 41.800 151.400 42.200 ;
        RECT 150.700 41.100 151.100 41.800 ;
        RECT 154.700 41.100 155.100 44.800 ;
        RECT 155.500 44.200 155.800 44.800 ;
        RECT 155.400 43.800 155.800 44.200 ;
        RECT 156.600 41.100 157.000 45.400 ;
        RECT 159.900 45.200 160.200 45.800 ;
        RECT 163.000 45.500 165.800 45.600 ;
        RECT 162.900 45.400 165.800 45.500 ;
        RECT 159.000 44.900 160.200 45.200 ;
        RECT 160.900 45.300 165.800 45.400 ;
        RECT 160.900 45.100 163.300 45.300 ;
        RECT 159.000 44.400 159.300 44.900 ;
        RECT 158.600 44.000 159.300 44.400 ;
        RECT 160.100 44.500 160.500 44.600 ;
        RECT 160.900 44.500 161.200 45.100 ;
        RECT 160.100 44.200 161.200 44.500 ;
        RECT 161.500 44.500 164.200 44.800 ;
        RECT 161.500 44.400 161.900 44.500 ;
        RECT 163.800 44.400 164.200 44.500 ;
        RECT 160.700 43.700 161.100 43.800 ;
        RECT 162.100 43.700 162.500 43.800 ;
        RECT 159.000 43.100 159.400 43.500 ;
        RECT 160.700 43.400 162.500 43.700 ;
        RECT 161.100 43.100 161.400 43.400 ;
        RECT 163.800 43.100 164.200 43.500 ;
        RECT 158.700 41.100 159.300 43.100 ;
        RECT 161.000 41.100 161.400 43.100 ;
        RECT 163.200 42.800 164.200 43.100 ;
        RECT 163.200 41.100 163.600 42.800 ;
        RECT 165.400 41.100 165.800 45.300 ;
        RECT 167.700 45.100 168.000 46.800 ;
        RECT 168.600 45.100 169.000 45.200 ;
        RECT 167.500 44.800 168.000 45.100 ;
        RECT 168.300 44.800 169.000 45.100 ;
        RECT 167.500 41.100 167.900 44.800 ;
        RECT 168.300 44.200 168.600 44.800 ;
        RECT 168.200 43.800 168.600 44.200 ;
        RECT 169.400 41.100 169.800 49.900 ;
        RECT 170.200 47.800 170.600 48.600 ;
        RECT 171.000 47.700 171.400 49.900 ;
        RECT 173.100 49.200 173.700 49.900 ;
        RECT 173.100 48.900 173.800 49.200 ;
        RECT 175.400 48.900 175.800 49.900 ;
        RECT 177.600 49.200 178.000 49.900 ;
        RECT 177.600 48.900 178.600 49.200 ;
        RECT 173.400 48.500 173.800 48.900 ;
        RECT 175.500 48.600 175.800 48.900 ;
        RECT 175.500 48.300 176.900 48.600 ;
        RECT 176.500 48.200 176.900 48.300 ;
        RECT 177.400 48.200 177.800 48.600 ;
        RECT 178.200 48.500 178.600 48.900 ;
        RECT 172.500 47.700 172.900 47.800 ;
        RECT 171.000 47.400 172.900 47.700 ;
        RECT 171.000 45.700 171.400 47.400 ;
        RECT 174.500 47.100 174.900 47.200 ;
        RECT 177.400 47.100 177.700 48.200 ;
        RECT 179.800 47.500 180.200 49.900 ;
        RECT 179.000 47.100 179.800 47.200 ;
        RECT 174.300 46.800 179.800 47.100 ;
        RECT 173.400 46.400 173.800 46.500 ;
        RECT 171.900 46.100 173.800 46.400 ;
        RECT 174.300 46.200 174.600 46.800 ;
        RECT 177.900 46.700 178.300 46.800 ;
        RECT 178.700 46.200 179.100 46.300 ;
        RECT 171.900 46.000 172.300 46.100 ;
        RECT 174.200 45.800 174.600 46.200 ;
        RECT 176.600 45.900 179.100 46.200 ;
        RECT 176.600 45.800 177.000 45.900 ;
        RECT 172.700 45.700 173.100 45.800 ;
        RECT 171.000 45.400 173.100 45.700 ;
        RECT 171.000 41.100 171.400 45.400 ;
        RECT 174.300 45.200 174.600 45.800 ;
        RECT 177.400 45.500 180.200 45.600 ;
        RECT 177.300 45.400 180.200 45.500 ;
        RECT 173.400 44.900 174.600 45.200 ;
        RECT 175.300 45.300 180.200 45.400 ;
        RECT 175.300 45.100 177.700 45.300 ;
        RECT 173.400 44.400 173.700 44.900 ;
        RECT 173.000 44.000 173.700 44.400 ;
        RECT 174.500 44.500 174.900 44.600 ;
        RECT 175.300 44.500 175.600 45.100 ;
        RECT 174.500 44.200 175.600 44.500 ;
        RECT 175.900 44.500 178.600 44.800 ;
        RECT 175.900 44.400 176.300 44.500 ;
        RECT 178.200 44.400 178.600 44.500 ;
        RECT 175.100 43.700 175.500 43.800 ;
        RECT 176.500 43.700 176.900 43.800 ;
        RECT 173.400 43.100 173.800 43.500 ;
        RECT 175.100 43.400 176.900 43.700 ;
        RECT 175.500 43.100 175.800 43.400 ;
        RECT 178.200 43.100 178.600 43.500 ;
        RECT 173.100 41.100 173.700 43.100 ;
        RECT 175.400 41.100 175.800 43.100 ;
        RECT 177.600 42.800 178.600 43.100 ;
        RECT 177.600 41.100 178.000 42.800 ;
        RECT 179.800 41.100 180.200 45.300 ;
        RECT 0.600 35.700 1.000 39.900 ;
        RECT 2.800 38.200 3.200 39.900 ;
        RECT 2.200 37.900 3.200 38.200 ;
        RECT 5.000 37.900 5.400 39.900 ;
        RECT 7.100 37.900 7.700 39.900 ;
        RECT 2.200 37.500 2.600 37.900 ;
        RECT 5.000 37.600 5.300 37.900 ;
        RECT 3.900 37.300 5.700 37.600 ;
        RECT 7.000 37.500 7.400 37.900 ;
        RECT 3.900 37.200 4.300 37.300 ;
        RECT 5.300 37.200 5.700 37.300 ;
        RECT 2.200 36.500 2.600 36.600 ;
        RECT 4.500 36.500 4.900 36.600 ;
        RECT 2.200 36.200 4.900 36.500 ;
        RECT 5.200 36.500 6.300 36.800 ;
        RECT 5.200 35.900 5.500 36.500 ;
        RECT 5.900 36.400 6.300 36.500 ;
        RECT 7.100 36.600 7.800 37.000 ;
        RECT 7.100 36.100 7.400 36.600 ;
        RECT 3.100 35.700 5.500 35.900 ;
        RECT 0.600 35.600 5.500 35.700 ;
        RECT 6.200 35.800 7.400 36.100 ;
        RECT 0.600 35.500 3.500 35.600 ;
        RECT 0.600 35.400 3.400 35.500 ;
        RECT 3.800 35.100 4.200 35.200 ;
        RECT 1.700 34.800 4.200 35.100 ;
        RECT 1.700 34.700 2.100 34.800 ;
        RECT 2.500 34.200 2.900 34.300 ;
        RECT 6.200 34.200 6.500 35.800 ;
        RECT 9.400 35.600 9.800 39.900 ;
        RECT 12.100 36.400 12.500 39.900 ;
        RECT 14.200 37.500 14.600 39.500 ;
        RECT 11.700 36.100 12.500 36.400 ;
        RECT 7.700 35.300 9.800 35.600 ;
        RECT 7.700 35.200 8.100 35.300 ;
        RECT 8.500 34.900 8.900 35.000 ;
        RECT 7.000 34.600 8.900 34.900 ;
        RECT 7.000 34.500 7.400 34.600 ;
        RECT 1.000 33.900 6.500 34.200 ;
        RECT 1.000 33.800 1.800 33.900 ;
        RECT 0.600 31.100 1.000 33.500 ;
        RECT 3.100 33.200 3.400 33.900 ;
        RECT 5.900 33.800 6.300 33.900 ;
        RECT 9.400 33.600 9.800 35.300 ;
        RECT 11.000 34.800 11.400 35.600 ;
        RECT 11.700 34.200 12.000 36.100 ;
        RECT 14.300 35.800 14.600 37.500 ;
        RECT 15.000 36.200 15.400 39.900 ;
        RECT 16.600 39.600 18.600 39.900 ;
        RECT 16.600 36.200 17.000 39.600 ;
        RECT 15.000 35.900 17.000 36.200 ;
        RECT 17.400 35.900 17.800 39.300 ;
        RECT 18.200 35.900 18.600 39.600 ;
        RECT 12.700 35.500 14.600 35.800 ;
        RECT 17.400 35.600 17.700 35.900 ;
        RECT 19.000 35.700 19.400 39.900 ;
        RECT 21.200 38.200 21.600 39.900 ;
        RECT 20.600 37.900 21.600 38.200 ;
        RECT 23.400 37.900 23.800 39.900 ;
        RECT 25.500 37.900 26.100 39.900 ;
        RECT 20.600 37.500 21.000 37.900 ;
        RECT 23.400 37.600 23.700 37.900 ;
        RECT 22.300 37.300 24.100 37.600 ;
        RECT 25.400 37.500 25.800 37.900 ;
        RECT 22.300 37.200 22.700 37.300 ;
        RECT 23.700 37.200 24.100 37.300 ;
        RECT 20.600 36.500 21.000 36.600 ;
        RECT 22.900 36.500 23.300 36.600 ;
        RECT 20.600 36.200 23.300 36.500 ;
        RECT 23.600 36.500 24.700 36.800 ;
        RECT 23.600 35.900 23.900 36.500 ;
        RECT 24.300 36.400 24.700 36.500 ;
        RECT 25.500 36.600 26.200 37.000 ;
        RECT 25.500 36.100 25.800 36.600 ;
        RECT 21.500 35.700 23.900 35.900 ;
        RECT 19.000 35.600 23.900 35.700 ;
        RECT 24.600 35.800 25.800 36.100 ;
        RECT 12.700 34.500 13.000 35.500 ;
        RECT 15.400 35.200 15.800 35.400 ;
        RECT 16.700 35.300 17.700 35.600 ;
        RECT 16.700 35.200 17.000 35.300 ;
        RECT 10.200 34.100 10.600 34.200 ;
        RECT 11.000 34.100 12.000 34.200 ;
        RECT 12.300 34.100 13.000 34.500 ;
        RECT 13.400 34.400 13.800 35.200 ;
        RECT 14.200 34.400 14.600 35.200 ;
        RECT 15.000 34.900 15.800 35.200 ;
        RECT 15.000 34.800 15.400 34.900 ;
        RECT 16.600 34.800 17.000 35.200 ;
        RECT 18.200 34.800 18.600 35.600 ;
        RECT 19.000 35.500 21.900 35.600 ;
        RECT 19.000 35.400 21.800 35.500 ;
        RECT 22.200 35.100 22.600 35.200 ;
        RECT 20.100 34.800 22.600 35.100 ;
        RECT 10.200 33.800 12.000 34.100 ;
        RECT 7.900 33.300 9.800 33.600 ;
        RECT 7.900 33.200 8.300 33.300 ;
        RECT 2.200 32.100 2.600 32.500 ;
        RECT 3.000 32.400 3.400 33.200 ;
        RECT 3.900 32.700 4.300 32.800 ;
        RECT 3.900 32.400 5.300 32.700 ;
        RECT 5.000 32.100 5.300 32.400 ;
        RECT 7.000 32.100 7.400 32.500 ;
        RECT 2.200 31.800 3.200 32.100 ;
        RECT 2.800 31.100 3.200 31.800 ;
        RECT 5.000 31.100 5.400 32.100 ;
        RECT 7.000 31.800 7.700 32.100 ;
        RECT 7.100 31.100 7.700 31.800 ;
        RECT 9.400 31.100 9.800 33.300 ;
        RECT 11.700 33.500 12.000 33.800 ;
        RECT 12.500 33.900 13.000 34.100 ;
        RECT 12.500 33.600 14.600 33.900 ;
        RECT 15.800 33.800 16.200 34.600 ;
        RECT 11.700 33.300 12.100 33.500 ;
        RECT 11.700 33.000 12.500 33.300 ;
        RECT 12.100 31.500 12.500 33.000 ;
        RECT 14.300 32.500 14.600 33.600 ;
        RECT 16.700 33.100 17.000 34.800 ;
        RECT 17.300 34.400 17.700 34.800 ;
        RECT 20.100 34.700 20.500 34.800 ;
        RECT 17.400 34.200 17.700 34.400 ;
        RECT 20.900 34.200 21.300 34.300 ;
        RECT 24.600 34.200 24.900 35.800 ;
        RECT 27.800 35.600 28.200 39.900 ;
        RECT 26.100 35.300 28.200 35.600 ;
        RECT 28.600 37.500 29.000 39.500 ;
        RECT 28.600 35.800 28.900 37.500 ;
        RECT 30.700 36.400 31.100 39.900 ;
        RECT 30.700 36.100 31.500 36.400 ;
        RECT 28.600 35.500 30.500 35.800 ;
        RECT 26.100 35.200 26.500 35.300 ;
        RECT 26.900 34.900 27.300 35.000 ;
        RECT 25.400 34.600 27.300 34.900 ;
        RECT 25.400 34.500 25.800 34.600 ;
        RECT 17.400 33.800 17.800 34.200 ;
        RECT 19.400 33.900 24.900 34.200 ;
        RECT 19.400 33.800 20.200 33.900 ;
        RECT 14.200 31.500 14.600 32.500 ;
        RECT 16.500 31.100 17.300 33.100 ;
        RECT 19.000 31.100 19.400 33.500 ;
        RECT 21.500 33.200 21.800 33.900 ;
        RECT 24.300 33.800 24.700 33.900 ;
        RECT 27.800 33.600 28.200 35.300 ;
        RECT 28.600 34.400 29.000 35.200 ;
        RECT 29.400 34.400 29.800 35.200 ;
        RECT 30.200 34.500 30.500 35.500 ;
        RECT 30.200 34.100 30.900 34.500 ;
        RECT 31.200 34.200 31.500 36.100 ;
        RECT 31.800 35.100 32.200 35.600 ;
        RECT 33.400 35.100 33.800 39.900 ;
        RECT 35.000 37.500 35.400 39.500 ;
        RECT 35.000 35.800 35.300 37.500 ;
        RECT 37.100 36.400 37.500 39.900 ;
        RECT 37.100 36.100 37.900 36.400 ;
        RECT 35.000 35.500 36.900 35.800 ;
        RECT 31.800 34.800 33.800 35.100 ;
        RECT 30.200 33.900 30.700 34.100 ;
        RECT 26.300 33.300 28.200 33.600 ;
        RECT 26.300 33.200 26.700 33.300 ;
        RECT 20.600 32.100 21.000 32.500 ;
        RECT 21.400 32.400 21.800 33.200 ;
        RECT 22.300 32.700 22.700 32.800 ;
        RECT 22.300 32.400 23.700 32.700 ;
        RECT 23.400 32.100 23.700 32.400 ;
        RECT 25.400 32.100 25.800 32.500 ;
        RECT 20.600 31.800 21.600 32.100 ;
        RECT 21.200 31.100 21.600 31.800 ;
        RECT 23.400 31.100 23.800 32.100 ;
        RECT 25.400 31.800 26.100 32.100 ;
        RECT 25.500 31.100 26.100 31.800 ;
        RECT 27.800 31.100 28.200 33.300 ;
        RECT 28.600 33.600 30.700 33.900 ;
        RECT 31.200 33.800 32.200 34.200 ;
        RECT 28.600 32.500 28.900 33.600 ;
        RECT 31.200 33.500 31.500 33.800 ;
        RECT 31.100 33.300 31.500 33.500 ;
        RECT 30.700 33.200 31.500 33.300 ;
        RECT 30.200 33.000 31.500 33.200 ;
        RECT 30.200 32.800 31.100 33.000 ;
        RECT 28.600 31.500 29.000 32.500 ;
        RECT 30.700 31.500 31.100 32.800 ;
        RECT 33.400 31.100 33.800 34.800 ;
        RECT 35.000 34.400 35.400 35.200 ;
        RECT 35.800 34.400 36.200 35.200 ;
        RECT 36.600 34.500 36.900 35.500 ;
        RECT 36.600 34.100 37.300 34.500 ;
        RECT 37.600 34.200 37.900 36.100 ;
        RECT 38.200 35.100 38.600 35.600 ;
        RECT 41.400 35.100 41.800 39.900 ;
        RECT 43.000 37.900 43.400 39.900 ;
        RECT 43.100 37.800 43.400 37.900 ;
        RECT 44.600 37.900 45.000 39.900 ;
        RECT 44.600 37.800 44.900 37.900 ;
        RECT 43.100 37.500 44.900 37.800 ;
        RECT 47.000 37.800 47.400 39.900 ;
        RECT 48.600 37.900 49.000 39.900 ;
        RECT 50.200 37.900 50.600 39.900 ;
        RECT 48.600 37.800 48.900 37.900 ;
        RECT 47.000 37.500 48.900 37.800 ;
        RECT 50.300 37.800 50.600 37.900 ;
        RECT 51.800 37.900 52.200 39.900 ;
        RECT 51.800 37.800 52.100 37.900 ;
        RECT 50.300 37.500 52.100 37.800 ;
        RECT 43.100 36.200 43.400 37.500 ;
        RECT 43.800 36.400 44.200 37.200 ;
        RECT 47.000 37.100 47.300 37.500 ;
        RECT 45.400 36.800 47.300 37.100 ;
        RECT 43.000 35.800 43.400 36.200 ;
        RECT 38.200 34.800 41.800 35.100 ;
        RECT 36.600 33.900 37.100 34.100 ;
        RECT 35.000 33.600 37.100 33.900 ;
        RECT 37.600 33.800 38.600 34.200 ;
        RECT 34.200 32.400 34.600 33.200 ;
        RECT 35.000 32.500 35.300 33.600 ;
        RECT 37.600 33.500 37.900 33.800 ;
        RECT 37.500 33.300 37.900 33.500 ;
        RECT 37.100 33.000 37.900 33.300 ;
        RECT 35.000 31.500 35.400 32.500 ;
        RECT 37.100 32.200 37.500 33.000 ;
        RECT 37.100 31.800 37.800 32.200 ;
        RECT 37.100 31.500 37.500 31.800 ;
        RECT 41.400 31.100 41.800 34.800 ;
        RECT 43.100 34.200 43.400 35.800 ;
        RECT 45.400 36.200 45.700 36.800 ;
        RECT 47.800 36.400 48.200 37.200 ;
        RECT 48.600 36.200 48.900 37.500 ;
        RECT 51.000 36.400 51.400 37.200 ;
        RECT 51.800 36.200 52.100 37.500 ;
        RECT 45.400 35.400 45.800 36.200 ;
        RECT 46.200 35.400 46.600 36.200 ;
        RECT 48.600 35.800 49.000 36.200 ;
        RECT 44.200 34.800 45.000 35.200 ;
        RECT 47.000 34.800 47.800 35.200 ;
        RECT 48.600 34.200 48.900 35.800 ;
        RECT 49.400 34.800 49.800 36.200 ;
        RECT 51.800 35.800 52.200 36.200 ;
        RECT 50.200 34.800 51.000 35.200 ;
        RECT 51.800 34.200 52.100 35.800 ;
        RECT 43.100 34.100 43.900 34.200 ;
        RECT 48.100 34.100 48.900 34.200 ;
        RECT 51.300 34.100 52.100 34.200 ;
        RECT 43.100 33.900 44.000 34.100 ;
        RECT 42.200 32.400 42.600 33.200 ;
        RECT 43.600 31.100 44.000 33.900 ;
        RECT 48.000 33.900 48.900 34.100 ;
        RECT 51.200 33.900 52.100 34.100 ;
        RECT 48.000 31.100 48.400 33.900 ;
        RECT 51.200 31.100 51.600 33.900 ;
        RECT 52.600 31.100 53.000 39.900 ;
        RECT 55.000 37.900 55.400 39.900 ;
        RECT 55.100 37.800 55.400 37.900 ;
        RECT 56.600 37.900 57.000 39.900 ;
        RECT 56.600 37.800 56.900 37.900 ;
        RECT 55.100 37.500 56.900 37.800 ;
        RECT 55.800 36.400 56.200 37.200 ;
        RECT 56.600 36.200 56.900 37.500 ;
        RECT 57.700 36.300 58.100 39.900 ;
        RECT 60.100 39.200 60.500 39.900 ;
        RECT 59.800 38.800 60.500 39.200 ;
        RECT 54.200 35.400 54.600 36.200 ;
        RECT 56.600 35.800 57.000 36.200 ;
        RECT 57.700 35.900 58.600 36.300 ;
        RECT 60.100 36.200 60.500 38.800 ;
        RECT 59.800 35.900 60.500 36.200 ;
        RECT 55.000 34.800 55.800 35.200 ;
        RECT 56.600 34.200 56.900 35.800 ;
        RECT 57.400 34.800 57.800 35.600 ;
        RECT 58.200 35.100 58.500 35.900 ;
        RECT 59.800 35.200 60.100 35.900 ;
        RECT 62.200 35.600 62.600 39.900 ;
        RECT 60.600 35.400 62.600 35.600 ;
        RECT 60.500 35.300 62.600 35.400 ;
        RECT 63.800 36.100 64.200 39.900 ;
        RECT 64.600 36.800 65.000 37.200 ;
        RECT 64.600 36.100 64.900 36.800 ;
        RECT 63.800 35.800 64.900 36.100 ;
        RECT 59.000 35.100 59.400 35.200 ;
        RECT 58.200 34.800 59.400 35.100 ;
        RECT 59.800 34.800 60.200 35.200 ;
        RECT 60.500 35.000 60.900 35.300 ;
        RECT 53.400 33.400 53.800 34.200 ;
        RECT 56.100 34.100 56.900 34.200 ;
        RECT 56.000 33.900 56.900 34.100 ;
        RECT 58.200 34.200 58.500 34.800 ;
        RECT 56.000 31.100 56.400 33.900 ;
        RECT 58.200 33.800 58.600 34.200 ;
        RECT 58.200 32.100 58.500 33.800 ;
        RECT 59.000 32.400 59.400 33.200 ;
        RECT 59.800 33.100 60.100 34.800 ;
        RECT 60.500 33.500 60.800 35.000 ;
        RECT 60.500 33.200 61.700 33.500 ;
        RECT 58.200 31.100 58.600 32.100 ;
        RECT 59.800 31.100 60.200 33.100 ;
        RECT 61.400 32.100 61.700 33.200 ;
        RECT 61.400 31.100 61.800 32.100 ;
        RECT 63.800 31.100 64.200 35.800 ;
        RECT 65.400 33.100 65.800 39.900 ;
        RECT 67.000 36.900 67.400 39.900 ;
        RECT 67.100 36.600 67.400 36.900 ;
        RECT 68.600 39.600 70.600 39.900 ;
        RECT 68.600 36.900 69.000 39.600 ;
        RECT 69.400 36.900 69.800 39.300 ;
        RECT 70.200 37.000 70.600 39.600 ;
        RECT 71.100 39.600 72.900 39.900 ;
        RECT 71.100 39.500 71.400 39.600 ;
        RECT 68.600 36.600 68.900 36.900 ;
        RECT 66.200 35.800 66.600 36.600 ;
        RECT 67.100 36.300 68.900 36.600 ;
        RECT 69.500 36.700 69.800 36.900 ;
        RECT 71.000 36.700 71.400 39.500 ;
        RECT 72.600 39.500 72.900 39.600 ;
        RECT 69.500 36.500 71.400 36.700 ;
        RECT 71.800 36.500 72.200 39.300 ;
        RECT 72.600 36.500 73.000 39.500 ;
        RECT 69.500 36.400 71.300 36.500 ;
        RECT 71.800 36.200 72.100 36.500 ;
        RECT 71.800 36.100 72.200 36.200 ;
        RECT 70.500 35.800 72.200 36.100 ;
        RECT 69.400 34.800 70.200 35.200 ;
        RECT 65.400 32.800 66.300 33.100 ;
        RECT 67.800 32.800 68.700 33.200 ;
        RECT 65.900 31.100 66.300 32.800 ;
        RECT 70.500 32.500 70.800 35.800 ;
        RECT 72.600 35.100 73.000 35.200 ;
        RECT 74.200 35.100 74.600 39.900 ;
        RECT 76.100 36.300 76.500 39.900 ;
        RECT 79.500 38.200 79.900 39.900 ;
        RECT 80.900 39.200 81.300 39.900 ;
        RECT 83.000 39.600 85.000 39.900 ;
        RECT 80.900 38.800 81.800 39.200 ;
        RECT 79.500 37.800 80.200 38.200 ;
        RECT 79.500 36.300 79.900 37.800 ;
        RECT 76.100 35.900 77.000 36.300 ;
        RECT 79.000 35.900 79.900 36.300 ;
        RECT 80.900 36.300 81.300 38.800 ;
        RECT 80.900 35.900 81.800 36.300 ;
        RECT 83.000 35.900 83.400 39.600 ;
        RECT 83.800 35.900 84.200 39.300 ;
        RECT 84.600 36.200 85.000 39.600 ;
        RECT 86.200 36.200 86.600 39.900 ;
        RECT 84.600 35.900 86.600 36.200 ;
        RECT 88.600 37.500 89.000 39.500 ;
        RECT 72.600 34.800 74.600 35.100 ;
        RECT 75.800 34.800 76.200 35.600 ;
        RECT 76.600 35.100 76.900 35.900 ;
        RECT 76.600 34.800 77.700 35.100 ;
        RECT 74.200 33.100 74.600 34.800 ;
        RECT 68.800 32.200 70.800 32.500 ;
        RECT 68.800 32.100 69.100 32.200 ;
        RECT 68.600 31.800 69.100 32.100 ;
        RECT 70.200 32.100 70.800 32.200 ;
        RECT 73.700 32.800 74.600 33.100 ;
        RECT 76.600 34.200 76.900 34.800 ;
        RECT 77.400 34.200 77.700 34.800 ;
        RECT 79.100 34.200 79.400 35.900 ;
        RECT 79.800 34.800 80.200 35.600 ;
        RECT 80.600 34.800 81.000 35.600 ;
        RECT 76.600 33.800 77.000 34.200 ;
        RECT 77.400 33.800 77.800 34.200 ;
        RECT 79.000 33.800 79.400 34.200 ;
        RECT 68.600 31.100 69.000 31.800 ;
        RECT 70.200 31.100 70.600 32.100 ;
        RECT 73.700 31.100 74.100 32.800 ;
        RECT 76.600 32.100 76.900 33.800 ;
        RECT 77.400 33.100 77.800 33.200 ;
        RECT 78.200 33.100 78.600 33.200 ;
        RECT 77.400 32.800 78.600 33.100 ;
        RECT 77.400 32.400 77.800 32.800 ;
        RECT 78.200 32.400 78.600 32.800 ;
        RECT 79.100 32.200 79.400 33.800 ;
        RECT 76.600 31.100 77.000 32.100 ;
        RECT 79.000 31.100 79.400 32.200 ;
        RECT 81.400 34.200 81.700 35.900 ;
        RECT 83.900 35.600 84.200 35.900 ;
        RECT 88.600 35.800 88.900 37.500 ;
        RECT 90.700 36.400 91.100 39.900 ;
        RECT 90.700 36.100 91.500 36.400 ;
        RECT 91.000 35.800 91.500 36.100 ;
        RECT 83.000 34.800 83.400 35.600 ;
        RECT 83.900 35.300 84.900 35.600 ;
        RECT 88.600 35.500 90.500 35.800 ;
        RECT 84.600 35.200 84.900 35.300 ;
        RECT 85.800 35.200 86.200 35.400 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 85.800 35.100 86.600 35.200 ;
        RECT 87.000 35.100 87.400 35.200 ;
        RECT 85.800 34.900 87.400 35.100 ;
        RECT 86.200 34.800 87.400 34.900 ;
        RECT 83.900 34.400 84.300 34.800 ;
        RECT 83.900 34.200 84.200 34.400 ;
        RECT 81.400 33.800 81.800 34.200 ;
        RECT 83.800 33.800 84.200 34.200 ;
        RECT 81.400 32.100 81.700 33.800 ;
        RECT 82.200 32.400 82.600 33.200 ;
        RECT 84.600 33.100 84.900 34.800 ;
        RECT 85.400 33.800 85.800 34.600 ;
        RECT 88.600 34.400 89.000 35.200 ;
        RECT 89.400 34.400 89.800 35.200 ;
        RECT 90.200 34.500 90.500 35.500 ;
        RECT 90.200 34.100 90.900 34.500 ;
        RECT 91.200 34.200 91.500 35.800 ;
        RECT 91.800 35.100 92.200 35.600 ;
        RECT 93.400 35.100 93.800 39.900 ;
        RECT 95.000 35.700 95.400 39.900 ;
        RECT 97.200 38.200 97.600 39.900 ;
        RECT 96.600 37.900 97.600 38.200 ;
        RECT 99.400 37.900 99.800 39.900 ;
        RECT 101.500 37.900 102.100 39.900 ;
        RECT 96.600 37.500 97.000 37.900 ;
        RECT 99.400 37.600 99.700 37.900 ;
        RECT 98.300 37.300 100.100 37.600 ;
        RECT 101.400 37.500 101.800 37.900 ;
        RECT 98.300 37.200 98.700 37.300 ;
        RECT 99.700 37.200 100.100 37.300 ;
        RECT 96.600 36.500 97.000 36.600 ;
        RECT 98.900 36.500 99.300 36.600 ;
        RECT 96.600 36.200 99.300 36.500 ;
        RECT 99.600 36.500 100.700 36.800 ;
        RECT 99.600 35.900 99.900 36.500 ;
        RECT 100.300 36.400 100.700 36.500 ;
        RECT 101.500 36.600 102.200 37.000 ;
        RECT 101.500 36.100 101.800 36.600 ;
        RECT 97.500 35.700 99.900 35.900 ;
        RECT 95.000 35.600 99.900 35.700 ;
        RECT 100.600 35.800 101.800 36.100 ;
        RECT 95.000 35.500 97.900 35.600 ;
        RECT 95.000 35.400 97.800 35.500 ;
        RECT 98.200 35.100 98.600 35.200 ;
        RECT 91.800 34.800 93.800 35.100 ;
        RECT 90.200 33.900 90.700 34.100 ;
        RECT 88.600 33.600 90.700 33.900 ;
        RECT 91.200 33.800 92.200 34.200 ;
        RECT 81.400 31.100 81.800 32.100 ;
        RECT 84.300 31.100 85.100 33.100 ;
        RECT 88.600 32.500 88.900 33.600 ;
        RECT 91.200 33.500 91.500 33.800 ;
        RECT 91.100 33.300 91.500 33.500 ;
        RECT 90.700 33.000 91.500 33.300 ;
        RECT 88.600 31.500 89.000 32.500 ;
        RECT 90.700 31.500 91.100 33.000 ;
        RECT 93.400 31.100 93.800 34.800 ;
        RECT 96.100 34.800 98.600 35.100 ;
        RECT 96.100 34.700 96.500 34.800 ;
        RECT 97.400 34.700 97.800 34.800 ;
        RECT 96.900 34.200 97.300 34.300 ;
        RECT 100.600 34.200 100.900 35.800 ;
        RECT 103.800 35.600 104.200 39.900 ;
        RECT 105.900 36.300 106.300 39.900 ;
        RECT 105.400 35.900 106.300 36.300 ;
        RECT 107.000 35.900 107.400 39.900 ;
        RECT 107.800 36.200 108.200 39.900 ;
        RECT 109.400 36.200 109.800 39.900 ;
        RECT 107.800 35.900 109.800 36.200 ;
        RECT 102.100 35.300 104.200 35.600 ;
        RECT 102.100 35.200 102.500 35.300 ;
        RECT 102.900 34.900 103.300 35.000 ;
        RECT 101.400 34.600 103.300 34.900 ;
        RECT 101.400 34.500 101.800 34.600 ;
        RECT 95.400 33.900 100.900 34.200 ;
        RECT 95.400 33.800 96.200 33.900 ;
        RECT 94.200 32.400 94.600 33.200 ;
        RECT 95.000 31.100 95.400 33.500 ;
        RECT 97.500 32.800 97.800 33.900 ;
        RECT 100.300 33.800 100.700 33.900 ;
        RECT 103.800 33.600 104.200 35.300 ;
        RECT 105.500 34.200 105.800 35.900 ;
        RECT 106.200 34.800 106.600 35.600 ;
        RECT 107.100 35.200 107.400 35.900 ;
        RECT 110.200 35.600 110.600 39.900 ;
        RECT 112.300 37.900 112.900 39.900 ;
        RECT 114.600 37.900 115.000 39.900 ;
        RECT 116.800 38.200 117.200 39.900 ;
        RECT 116.800 37.900 117.800 38.200 ;
        RECT 112.600 37.500 113.000 37.900 ;
        RECT 114.700 37.600 115.000 37.900 ;
        RECT 114.300 37.300 116.100 37.600 ;
        RECT 117.400 37.500 117.800 37.900 ;
        RECT 114.300 37.200 114.700 37.300 ;
        RECT 115.700 37.200 116.100 37.300 ;
        RECT 112.200 36.600 112.900 37.000 ;
        RECT 112.600 36.100 112.900 36.600 ;
        RECT 113.700 36.500 114.800 36.800 ;
        RECT 113.700 36.400 114.100 36.500 ;
        RECT 112.600 35.800 113.800 36.100 ;
        RECT 109.000 35.200 109.400 35.400 ;
        RECT 110.200 35.300 112.300 35.600 ;
        RECT 107.000 34.900 108.200 35.200 ;
        RECT 109.000 34.900 109.800 35.200 ;
        RECT 107.000 34.800 107.400 34.900 ;
        RECT 105.400 33.800 105.800 34.200 ;
        RECT 102.300 33.300 104.200 33.600 ;
        RECT 102.300 33.200 102.700 33.300 ;
        RECT 96.600 32.100 97.000 32.500 ;
        RECT 97.400 32.400 97.800 32.800 ;
        RECT 98.300 32.700 98.700 32.800 ;
        RECT 98.300 32.400 99.700 32.700 ;
        RECT 99.400 32.100 99.700 32.400 ;
        RECT 101.400 32.100 101.800 32.500 ;
        RECT 96.600 31.800 97.600 32.100 ;
        RECT 97.200 31.100 97.600 31.800 ;
        RECT 99.400 31.100 99.800 32.100 ;
        RECT 101.400 31.800 102.100 32.100 ;
        RECT 101.500 31.100 102.100 31.800 ;
        RECT 103.800 31.100 104.200 33.300 ;
        RECT 104.600 32.400 105.000 33.200 ;
        RECT 105.500 33.100 105.800 33.800 ;
        RECT 107.900 33.200 108.200 34.900 ;
        RECT 109.400 34.800 109.800 34.900 ;
        RECT 108.600 33.800 109.000 34.600 ;
        RECT 107.000 33.100 107.400 33.200 ;
        RECT 105.400 32.800 107.400 33.100 ;
        RECT 105.500 32.100 105.800 32.800 ;
        RECT 107.100 32.400 107.500 32.800 ;
        RECT 105.400 31.100 105.800 32.100 ;
        RECT 107.800 31.100 108.200 33.200 ;
        RECT 110.200 33.600 110.600 35.300 ;
        RECT 111.900 35.200 112.300 35.300 ;
        RECT 111.100 34.900 111.500 35.000 ;
        RECT 111.100 34.600 113.000 34.900 ;
        RECT 112.600 34.500 113.000 34.600 ;
        RECT 113.500 34.200 113.800 35.800 ;
        RECT 114.500 35.900 114.800 36.500 ;
        RECT 115.100 36.500 115.500 36.600 ;
        RECT 117.400 36.500 117.800 36.600 ;
        RECT 115.100 36.200 117.800 36.500 ;
        RECT 114.500 35.700 116.900 35.900 ;
        RECT 119.000 35.700 119.400 39.900 ;
        RECT 121.100 39.200 121.500 39.900 ;
        RECT 120.600 38.800 121.500 39.200 ;
        RECT 121.100 36.200 121.500 38.800 ;
        RECT 121.800 36.800 122.200 37.200 ;
        RECT 121.900 36.200 122.200 36.800 ;
        RECT 121.100 35.900 121.600 36.200 ;
        RECT 121.900 35.900 122.600 36.200 ;
        RECT 114.500 35.600 119.400 35.700 ;
        RECT 116.500 35.500 119.400 35.600 ;
        RECT 116.600 35.400 119.400 35.500 ;
        RECT 114.200 35.100 114.600 35.200 ;
        RECT 115.800 35.100 116.200 35.200 ;
        RECT 114.200 34.800 118.300 35.100 ;
        RECT 117.900 34.700 118.300 34.800 ;
        RECT 120.600 34.400 121.000 35.200 ;
        RECT 117.100 34.200 117.500 34.300 ;
        RECT 121.300 34.200 121.600 35.900 ;
        RECT 122.200 35.800 122.600 35.900 ;
        RECT 123.000 35.600 123.400 39.900 ;
        RECT 125.100 39.200 125.500 39.900 ;
        RECT 125.100 38.800 125.800 39.200 ;
        RECT 125.100 36.200 125.500 38.800 ;
        RECT 125.100 35.900 125.800 36.200 ;
        RECT 123.000 35.400 125.000 35.600 ;
        RECT 123.000 35.300 125.100 35.400 ;
        RECT 124.700 35.000 125.100 35.300 ;
        RECT 125.500 35.200 125.800 35.900 ;
        RECT 127.000 35.600 127.400 39.900 ;
        RECT 128.600 35.600 129.000 39.900 ;
        RECT 130.200 35.600 130.600 39.900 ;
        RECT 131.800 35.600 132.200 39.900 ;
        RECT 124.000 34.200 124.400 34.600 ;
        RECT 113.500 33.900 119.000 34.200 ;
        RECT 113.700 33.800 114.100 33.900 ;
        RECT 115.800 33.800 116.200 33.900 ;
        RECT 110.200 33.300 112.100 33.600 ;
        RECT 110.200 31.100 110.600 33.300 ;
        RECT 111.700 33.200 112.100 33.300 ;
        RECT 116.600 32.800 116.900 33.900 ;
        RECT 118.200 33.800 119.000 33.900 ;
        RECT 119.800 34.100 120.200 34.200 ;
        RECT 119.800 33.800 120.600 34.100 ;
        RECT 121.300 33.800 122.600 34.200 ;
        RECT 123.800 33.800 124.300 34.200 ;
        RECT 120.200 33.600 120.600 33.800 ;
        RECT 115.700 32.700 116.100 32.800 ;
        RECT 112.600 32.100 113.000 32.500 ;
        RECT 114.700 32.400 116.100 32.700 ;
        RECT 116.600 32.400 117.000 32.800 ;
        RECT 114.700 32.100 115.000 32.400 ;
        RECT 117.400 32.100 117.800 32.500 ;
        RECT 112.300 31.800 113.000 32.100 ;
        RECT 112.300 31.100 112.900 31.800 ;
        RECT 114.600 31.100 115.000 32.100 ;
        RECT 116.800 31.800 117.800 32.100 ;
        RECT 116.800 31.100 117.200 31.800 ;
        RECT 119.000 31.100 119.400 33.500 ;
        RECT 119.900 33.100 121.700 33.300 ;
        RECT 122.200 33.100 122.500 33.800 ;
        RECT 124.800 33.500 125.100 35.000 ;
        RECT 125.400 34.800 125.800 35.200 ;
        RECT 123.900 33.200 125.100 33.500 ;
        RECT 119.800 33.000 121.800 33.100 ;
        RECT 119.800 31.100 120.200 33.000 ;
        RECT 121.400 31.100 121.800 33.000 ;
        RECT 122.200 31.100 122.600 33.100 ;
        RECT 123.000 32.400 123.400 33.200 ;
        RECT 123.900 32.100 124.200 33.200 ;
        RECT 125.500 33.100 125.800 34.800 ;
        RECT 126.200 35.200 127.400 35.600 ;
        RECT 127.900 35.200 129.000 35.600 ;
        RECT 129.500 35.200 130.600 35.600 ;
        RECT 131.300 35.200 132.200 35.600 ;
        RECT 133.400 35.700 133.800 39.900 ;
        RECT 135.600 38.200 136.000 39.900 ;
        RECT 135.000 37.900 136.000 38.200 ;
        RECT 137.800 37.900 138.200 39.900 ;
        RECT 139.900 37.900 140.500 39.900 ;
        RECT 135.000 37.500 135.400 37.900 ;
        RECT 137.800 37.600 138.100 37.900 ;
        RECT 136.700 37.300 138.500 37.600 ;
        RECT 139.800 37.500 140.200 37.900 ;
        RECT 136.700 37.200 137.100 37.300 ;
        RECT 138.100 37.200 138.500 37.300 ;
        RECT 135.000 36.500 135.400 36.600 ;
        RECT 137.300 36.500 137.700 36.600 ;
        RECT 135.000 36.200 137.700 36.500 ;
        RECT 138.000 36.500 139.100 36.800 ;
        RECT 138.000 35.900 138.300 36.500 ;
        RECT 138.700 36.400 139.100 36.500 ;
        RECT 139.900 36.600 140.600 37.000 ;
        RECT 139.900 36.100 140.200 36.600 ;
        RECT 135.900 35.700 138.300 35.900 ;
        RECT 133.400 35.600 138.300 35.700 ;
        RECT 139.000 35.800 140.200 36.100 ;
        RECT 133.400 35.500 136.300 35.600 ;
        RECT 133.400 35.400 136.200 35.500 ;
        RECT 126.200 33.800 126.600 35.200 ;
        RECT 127.900 34.500 128.300 35.200 ;
        RECT 129.500 34.500 129.900 35.200 ;
        RECT 131.300 34.500 131.700 35.200 ;
        RECT 136.600 35.100 137.000 35.200 ;
        RECT 134.500 34.800 137.000 35.100 ;
        RECT 134.500 34.700 134.900 34.800 ;
        RECT 135.800 34.700 136.200 34.800 ;
        RECT 127.000 34.100 128.300 34.500 ;
        RECT 128.700 34.100 129.900 34.500 ;
        RECT 130.400 34.100 131.700 34.500 ;
        RECT 135.300 34.200 135.700 34.300 ;
        RECT 139.000 34.200 139.300 35.800 ;
        RECT 142.200 35.600 142.600 39.900 ;
        RECT 145.700 39.200 146.100 39.900 ;
        RECT 145.700 38.800 146.600 39.200 ;
        RECT 145.000 36.800 145.400 37.200 ;
        RECT 145.000 36.200 145.300 36.800 ;
        RECT 145.700 36.200 146.100 38.800 ;
        RECT 143.000 36.100 143.400 36.200 ;
        RECT 144.600 36.100 145.300 36.200 ;
        RECT 143.000 35.900 145.300 36.100 ;
        RECT 145.600 35.900 146.100 36.200 ;
        RECT 143.000 35.800 145.000 35.900 ;
        RECT 140.500 35.300 142.600 35.600 ;
        RECT 140.500 35.200 140.900 35.300 ;
        RECT 141.300 34.900 141.700 35.000 ;
        RECT 139.800 34.600 141.700 34.900 ;
        RECT 139.800 34.500 140.200 34.600 ;
        RECT 127.900 33.800 128.300 34.100 ;
        RECT 129.500 33.800 129.900 34.100 ;
        RECT 131.300 33.800 131.700 34.100 ;
        RECT 133.800 33.900 139.300 34.200 ;
        RECT 133.800 33.800 134.600 33.900 ;
        RECT 126.200 33.400 127.400 33.800 ;
        RECT 127.900 33.400 129.000 33.800 ;
        RECT 129.500 33.400 130.600 33.800 ;
        RECT 131.300 33.400 132.200 33.800 ;
        RECT 123.800 31.100 124.200 32.100 ;
        RECT 125.400 31.100 125.800 33.100 ;
        RECT 127.000 31.100 127.400 33.400 ;
        RECT 128.600 31.100 129.000 33.400 ;
        RECT 130.200 31.100 130.600 33.400 ;
        RECT 131.800 31.100 132.200 33.400 ;
        RECT 133.400 31.100 133.800 33.500 ;
        RECT 135.900 32.800 136.200 33.900 ;
        RECT 138.700 33.800 139.100 33.900 ;
        RECT 142.200 33.600 142.600 35.300 ;
        RECT 145.600 34.200 145.900 35.900 ;
        RECT 147.800 35.700 148.200 39.900 ;
        RECT 150.000 38.200 150.400 39.900 ;
        RECT 149.400 37.900 150.400 38.200 ;
        RECT 152.200 37.900 152.600 39.900 ;
        RECT 154.300 37.900 154.900 39.900 ;
        RECT 149.400 37.500 149.800 37.900 ;
        RECT 152.200 37.600 152.500 37.900 ;
        RECT 151.100 37.300 152.900 37.600 ;
        RECT 154.200 37.500 154.600 37.900 ;
        RECT 151.100 37.200 151.500 37.300 ;
        RECT 152.500 37.200 152.900 37.300 ;
        RECT 149.400 36.500 149.800 36.600 ;
        RECT 151.700 36.500 152.100 36.600 ;
        RECT 149.400 36.200 152.100 36.500 ;
        RECT 152.400 36.500 153.500 36.800 ;
        RECT 152.400 35.900 152.700 36.500 ;
        RECT 153.100 36.400 153.500 36.500 ;
        RECT 154.300 36.600 155.000 37.000 ;
        RECT 154.300 36.100 154.600 36.600 ;
        RECT 150.300 35.700 152.700 35.900 ;
        RECT 147.800 35.600 152.700 35.700 ;
        RECT 153.400 35.800 154.600 36.100 ;
        RECT 147.800 35.500 150.700 35.600 ;
        RECT 147.800 35.400 150.600 35.500 ;
        RECT 146.200 34.400 146.600 35.200 ;
        RECT 151.000 35.100 151.400 35.200 ;
        RECT 148.900 34.800 151.400 35.100 ;
        RECT 148.900 34.700 149.300 34.800 ;
        RECT 149.700 34.200 150.100 34.300 ;
        RECT 153.400 34.200 153.700 35.800 ;
        RECT 156.600 35.600 157.000 39.900 ;
        RECT 154.900 35.300 157.000 35.600 ;
        RECT 154.900 35.200 155.300 35.300 ;
        RECT 155.700 34.900 156.100 35.000 ;
        RECT 154.200 34.600 156.100 34.900 ;
        RECT 154.200 34.500 154.600 34.600 ;
        RECT 144.600 33.800 145.900 34.200 ;
        RECT 147.000 34.100 147.400 34.200 ;
        RECT 146.600 33.800 147.400 34.100 ;
        RECT 148.200 33.900 153.700 34.200 ;
        RECT 148.200 33.800 149.000 33.900 ;
        RECT 150.200 33.800 150.600 33.900 ;
        RECT 153.100 33.800 153.500 33.900 ;
        RECT 140.700 33.300 142.600 33.600 ;
        RECT 140.700 33.200 141.100 33.300 ;
        RECT 135.000 32.100 135.400 32.500 ;
        RECT 135.800 32.400 136.200 32.800 ;
        RECT 136.700 32.700 137.100 32.800 ;
        RECT 136.700 32.400 138.100 32.700 ;
        RECT 137.800 32.100 138.100 32.400 ;
        RECT 139.800 32.100 140.200 32.500 ;
        RECT 135.000 31.800 136.000 32.100 ;
        RECT 135.600 31.100 136.000 31.800 ;
        RECT 137.800 31.100 138.200 32.100 ;
        RECT 139.800 31.800 140.500 32.100 ;
        RECT 139.900 31.100 140.500 31.800 ;
        RECT 142.200 31.100 142.600 33.300 ;
        RECT 144.700 33.100 145.000 33.800 ;
        RECT 146.600 33.600 147.000 33.800 ;
        RECT 145.500 33.100 147.300 33.300 ;
        RECT 144.600 31.100 145.000 33.100 ;
        RECT 145.400 33.000 147.400 33.100 ;
        RECT 145.400 31.100 145.800 33.000 ;
        RECT 147.000 31.100 147.400 33.000 ;
        RECT 147.800 31.100 148.200 33.500 ;
        RECT 150.300 32.800 150.600 33.800 ;
        RECT 156.600 33.600 157.000 35.300 ;
        RECT 155.100 33.300 157.000 33.600 ;
        RECT 155.100 33.200 155.500 33.300 ;
        RECT 156.600 33.100 157.000 33.300 ;
        RECT 157.400 33.100 157.800 33.200 ;
        RECT 156.600 32.800 157.800 33.100 ;
        RECT 149.400 32.100 149.800 32.500 ;
        RECT 150.200 32.400 150.600 32.800 ;
        RECT 151.100 32.700 151.500 32.800 ;
        RECT 151.100 32.400 152.500 32.700 ;
        RECT 152.200 32.100 152.500 32.400 ;
        RECT 154.200 32.100 154.600 32.500 ;
        RECT 149.400 31.800 150.400 32.100 ;
        RECT 150.000 31.100 150.400 31.800 ;
        RECT 152.200 31.100 152.600 32.100 ;
        RECT 154.200 31.800 154.900 32.100 ;
        RECT 154.300 31.100 154.900 31.800 ;
        RECT 156.600 31.100 157.000 32.800 ;
        RECT 157.400 32.400 157.800 32.800 ;
        RECT 158.200 31.100 158.600 39.900 ;
        RECT 159.800 35.100 160.200 39.900 ;
        RECT 162.500 36.400 162.900 39.900 ;
        RECT 164.600 37.500 165.000 39.500 ;
        RECT 162.100 36.100 162.900 36.400 ;
        RECT 161.400 35.100 161.800 35.600 ;
        RECT 159.800 34.800 161.800 35.100 ;
        RECT 162.100 35.200 162.400 36.100 ;
        RECT 164.700 35.800 165.000 37.500 ;
        RECT 163.100 35.500 165.000 35.800 ;
        RECT 165.400 35.600 165.800 39.900 ;
        RECT 167.500 37.900 168.100 39.900 ;
        RECT 169.800 37.900 170.200 39.900 ;
        RECT 172.000 38.200 172.400 39.900 ;
        RECT 172.000 37.900 173.000 38.200 ;
        RECT 167.800 37.500 168.200 37.900 ;
        RECT 169.900 37.600 170.200 37.900 ;
        RECT 169.500 37.300 171.300 37.600 ;
        RECT 172.600 37.500 173.000 37.900 ;
        RECT 169.500 37.200 169.900 37.300 ;
        RECT 170.900 37.200 171.300 37.300 ;
        RECT 167.400 36.600 168.100 37.000 ;
        RECT 167.800 36.100 168.100 36.600 ;
        RECT 168.900 36.500 170.000 36.800 ;
        RECT 168.900 36.400 169.300 36.500 ;
        RECT 167.800 35.800 169.000 36.100 ;
        RECT 162.100 34.800 162.600 35.200 ;
        RECT 159.000 32.400 159.400 33.200 ;
        RECT 159.800 31.100 160.200 34.800 ;
        RECT 162.100 34.200 162.400 34.800 ;
        RECT 163.100 34.500 163.400 35.500 ;
        RECT 165.400 35.300 167.500 35.600 ;
        RECT 161.400 33.800 162.400 34.200 ;
        RECT 162.700 34.100 163.400 34.500 ;
        RECT 163.800 34.400 164.200 35.200 ;
        RECT 164.600 34.400 165.000 35.200 ;
        RECT 162.100 33.500 162.400 33.800 ;
        RECT 162.900 33.900 163.400 34.100 ;
        RECT 162.900 33.600 165.000 33.900 ;
        RECT 162.100 33.300 162.500 33.500 ;
        RECT 162.100 33.000 162.900 33.300 ;
        RECT 162.500 31.500 162.900 33.000 ;
        RECT 164.700 32.500 165.000 33.600 ;
        RECT 164.600 31.500 165.000 32.500 ;
        RECT 165.400 33.600 165.800 35.300 ;
        RECT 167.100 35.200 167.500 35.300 ;
        RECT 168.700 35.100 169.000 35.800 ;
        RECT 169.700 35.900 170.000 36.500 ;
        RECT 170.300 36.500 170.700 36.600 ;
        RECT 172.600 36.500 173.000 36.600 ;
        RECT 170.300 36.200 173.000 36.500 ;
        RECT 169.700 35.700 172.100 35.900 ;
        RECT 174.200 35.700 174.600 39.900 ;
        RECT 169.700 35.600 174.600 35.700 ;
        RECT 171.700 35.500 174.600 35.600 ;
        RECT 175.000 37.500 175.400 39.500 ;
        RECT 177.100 39.200 177.500 39.900 ;
        RECT 176.600 38.800 177.500 39.200 ;
        RECT 175.000 35.800 175.300 37.500 ;
        RECT 177.100 36.400 177.500 38.800 ;
        RECT 177.100 36.100 177.900 36.400 ;
        RECT 175.000 35.500 176.900 35.800 ;
        RECT 171.800 35.400 174.600 35.500 ;
        RECT 169.400 35.100 169.800 35.200 ;
        RECT 166.300 34.900 166.700 35.000 ;
        RECT 166.300 34.600 168.200 34.900 ;
        RECT 168.600 34.800 169.800 35.100 ;
        RECT 171.000 35.100 171.400 35.200 ;
        RECT 171.000 34.800 173.500 35.100 ;
        RECT 167.800 34.500 168.200 34.600 ;
        RECT 168.700 34.200 169.000 34.800 ;
        RECT 173.100 34.700 173.500 34.800 ;
        RECT 175.000 34.400 175.400 35.200 ;
        RECT 175.800 34.400 176.200 35.200 ;
        RECT 176.600 34.500 176.900 35.500 ;
        RECT 172.300 34.200 172.700 34.300 ;
        RECT 168.700 33.900 174.200 34.200 ;
        RECT 176.600 34.100 177.300 34.500 ;
        RECT 177.600 34.200 177.900 36.100 ;
        RECT 178.200 34.800 178.600 35.600 ;
        RECT 176.600 33.900 177.100 34.100 ;
        RECT 168.900 33.800 169.300 33.900 ;
        RECT 165.400 33.300 167.300 33.600 ;
        RECT 165.400 31.100 165.800 33.300 ;
        RECT 166.900 33.200 167.300 33.300 ;
        RECT 171.800 32.800 172.100 33.900 ;
        RECT 173.400 33.800 174.200 33.900 ;
        RECT 175.000 33.600 177.100 33.900 ;
        RECT 177.600 33.800 178.600 34.200 ;
        RECT 170.900 32.700 171.300 32.800 ;
        RECT 167.800 32.100 168.200 32.500 ;
        RECT 169.900 32.400 171.300 32.700 ;
        RECT 171.800 32.400 172.200 32.800 ;
        RECT 169.900 32.100 170.200 32.400 ;
        RECT 172.600 32.100 173.000 32.500 ;
        RECT 167.500 31.800 168.200 32.100 ;
        RECT 167.500 31.100 168.100 31.800 ;
        RECT 169.800 31.100 170.200 32.100 ;
        RECT 172.000 31.800 173.000 32.100 ;
        RECT 172.000 31.100 172.400 31.800 ;
        RECT 174.200 31.100 174.600 33.500 ;
        RECT 175.000 32.500 175.300 33.600 ;
        RECT 177.600 33.500 177.900 33.800 ;
        RECT 177.500 33.300 177.900 33.500 ;
        RECT 177.100 33.000 177.900 33.300 ;
        RECT 175.000 31.500 175.400 32.500 ;
        RECT 177.100 31.500 177.500 33.000 ;
        RECT 0.600 27.500 1.000 29.900 ;
        RECT 2.800 29.200 3.200 29.900 ;
        RECT 2.200 28.900 3.200 29.200 ;
        RECT 5.000 28.900 5.400 29.900 ;
        RECT 7.100 29.200 7.700 29.900 ;
        RECT 7.000 28.900 7.700 29.200 ;
        RECT 2.200 28.500 2.600 28.900 ;
        RECT 5.000 28.600 5.300 28.900 ;
        RECT 3.000 27.800 3.400 28.600 ;
        RECT 3.900 28.300 5.300 28.600 ;
        RECT 7.000 28.500 7.400 28.900 ;
        RECT 3.900 28.200 4.300 28.300 ;
        RECT 9.400 28.100 9.800 29.900 ;
        RECT 10.200 28.100 10.600 28.600 ;
        RECT 9.400 27.800 10.600 28.100 ;
        RECT 1.000 27.100 1.800 27.200 ;
        RECT 3.100 27.100 3.400 27.800 ;
        RECT 7.900 27.700 8.300 27.800 ;
        RECT 9.400 27.700 9.800 27.800 ;
        RECT 7.900 27.400 9.800 27.700 ;
        RECT 5.900 27.100 6.300 27.200 ;
        RECT 1.000 26.800 6.500 27.100 ;
        RECT 2.500 26.700 2.900 26.800 ;
        RECT 1.700 26.200 2.100 26.300 ;
        RECT 6.200 26.200 6.500 26.800 ;
        RECT 7.000 26.400 7.400 26.500 ;
        RECT 1.700 25.900 4.200 26.200 ;
        RECT 3.800 25.800 4.200 25.900 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 7.000 26.100 8.900 26.400 ;
        RECT 8.500 26.000 8.900 26.100 ;
        RECT 0.600 25.500 3.400 25.600 ;
        RECT 0.600 25.400 3.500 25.500 ;
        RECT 0.600 25.300 5.500 25.400 ;
        RECT 0.600 21.100 1.000 25.300 ;
        RECT 3.100 25.100 5.500 25.300 ;
        RECT 2.200 24.500 4.900 24.800 ;
        RECT 2.200 24.400 2.600 24.500 ;
        RECT 4.500 24.400 4.900 24.500 ;
        RECT 5.200 24.500 5.500 25.100 ;
        RECT 6.200 25.200 6.500 25.800 ;
        RECT 7.700 25.700 8.100 25.800 ;
        RECT 9.400 25.700 9.800 27.400 ;
        RECT 7.700 25.400 9.800 25.700 ;
        RECT 6.200 24.900 7.400 25.200 ;
        RECT 5.900 24.500 6.300 24.600 ;
        RECT 5.200 24.200 6.300 24.500 ;
        RECT 7.100 24.400 7.400 24.900 ;
        RECT 7.100 24.000 7.800 24.400 ;
        RECT 3.900 23.700 4.300 23.800 ;
        RECT 5.300 23.700 5.700 23.800 ;
        RECT 2.200 23.100 2.600 23.500 ;
        RECT 3.900 23.400 5.700 23.700 ;
        RECT 5.000 23.100 5.300 23.400 ;
        RECT 7.000 23.100 7.400 23.500 ;
        RECT 2.200 22.800 3.200 23.100 ;
        RECT 2.800 21.100 3.200 22.800 ;
        RECT 5.000 21.100 5.400 23.100 ;
        RECT 7.100 21.100 7.700 23.100 ;
        RECT 9.400 21.100 9.800 25.400 ;
        RECT 11.000 26.100 11.400 29.900 ;
        RECT 13.700 28.000 14.100 29.500 ;
        RECT 15.800 28.500 16.200 29.500 ;
        RECT 13.300 27.700 14.100 28.000 ;
        RECT 13.300 27.500 13.700 27.700 ;
        RECT 13.300 27.200 13.600 27.500 ;
        RECT 15.900 27.400 16.200 28.500 ;
        RECT 18.100 29.200 18.900 29.900 ;
        RECT 18.100 28.800 19.400 29.200 ;
        RECT 18.100 27.900 18.900 28.800 ;
        RECT 11.800 27.100 12.200 27.200 ;
        RECT 12.600 27.100 13.600 27.200 ;
        RECT 11.800 26.800 13.600 27.100 ;
        RECT 14.100 27.100 16.200 27.400 ;
        RECT 14.100 26.900 14.600 27.100 ;
        RECT 12.600 26.100 13.000 26.200 ;
        RECT 11.000 25.800 13.000 26.100 ;
        RECT 11.000 21.100 11.400 25.800 ;
        RECT 12.600 25.400 13.000 25.800 ;
        RECT 13.300 24.900 13.600 26.800 ;
        RECT 13.900 26.500 14.600 26.900 ;
        RECT 14.300 25.500 14.600 26.500 ;
        RECT 15.000 25.800 15.400 26.600 ;
        RECT 15.800 25.800 16.200 26.600 ;
        RECT 17.400 26.400 17.800 27.200 ;
        RECT 18.300 26.200 18.600 27.900 ;
        RECT 21.400 27.600 21.800 29.900 ;
        RECT 23.000 27.600 23.400 29.900 ;
        RECT 24.600 27.600 25.000 29.900 ;
        RECT 26.200 27.600 26.600 29.900 ;
        RECT 20.600 27.200 21.800 27.600 ;
        RECT 22.300 27.200 23.400 27.600 ;
        RECT 23.900 27.200 25.000 27.600 ;
        RECT 25.700 27.200 26.600 27.600 ;
        RECT 27.800 27.500 28.200 29.900 ;
        RECT 30.000 29.200 30.400 29.900 ;
        RECT 29.400 28.900 30.400 29.200 ;
        RECT 32.200 28.900 32.600 29.900 ;
        RECT 34.300 29.200 34.900 29.900 ;
        RECT 34.200 28.900 34.900 29.200 ;
        RECT 29.400 28.500 29.800 28.900 ;
        RECT 32.200 28.600 32.500 28.900 ;
        RECT 30.200 28.200 30.600 28.600 ;
        RECT 31.100 28.300 32.500 28.600 ;
        RECT 34.200 28.500 34.600 28.900 ;
        RECT 31.100 28.200 31.500 28.300 ;
        RECT 19.000 26.800 19.400 27.200 ;
        RECT 19.000 26.600 19.300 26.800 ;
        RECT 18.900 26.200 19.300 26.600 ;
        RECT 16.600 26.100 17.000 26.200 ;
        RECT 16.600 25.800 17.400 26.100 ;
        RECT 18.200 25.800 18.600 26.200 ;
        RECT 17.000 25.600 17.400 25.800 ;
        RECT 18.300 25.700 18.600 25.800 ;
        RECT 14.300 25.200 16.200 25.500 ;
        RECT 18.300 25.400 19.300 25.700 ;
        RECT 19.800 25.400 20.200 26.200 ;
        RECT 20.600 25.800 21.000 27.200 ;
        RECT 22.300 26.900 22.700 27.200 ;
        RECT 23.900 26.900 24.300 27.200 ;
        RECT 25.700 26.900 26.100 27.200 ;
        RECT 21.400 26.500 22.700 26.900 ;
        RECT 23.100 26.500 24.300 26.900 ;
        RECT 24.800 26.500 26.100 26.900 ;
        RECT 28.200 27.100 29.000 27.200 ;
        RECT 30.300 27.100 30.600 28.200 ;
        RECT 35.100 27.700 35.500 27.800 ;
        RECT 36.600 27.700 37.000 29.900 ;
        RECT 40.300 29.200 40.700 29.900 ;
        RECT 40.300 28.800 41.000 29.200 ;
        RECT 40.300 28.200 40.700 28.800 ;
        RECT 35.100 27.400 37.000 27.700 ;
        RECT 39.800 27.900 40.700 28.200 ;
        RECT 42.700 27.900 43.500 29.900 ;
        RECT 45.700 29.200 46.100 29.900 ;
        RECT 45.400 28.800 46.100 29.200 ;
        RECT 45.700 28.200 46.100 28.800 ;
        RECT 45.700 27.900 46.600 28.200 ;
        RECT 33.100 27.100 33.500 27.200 ;
        RECT 28.200 26.800 33.700 27.100 ;
        RECT 29.700 26.700 30.100 26.800 ;
        RECT 22.300 25.800 22.700 26.500 ;
        RECT 23.900 25.800 24.300 26.500 ;
        RECT 25.700 25.800 26.100 26.500 ;
        RECT 28.900 26.200 29.300 26.300 ;
        RECT 33.400 26.200 33.700 26.800 ;
        RECT 34.200 26.400 34.600 26.500 ;
        RECT 28.900 25.900 31.400 26.200 ;
        RECT 31.000 25.800 31.400 25.900 ;
        RECT 33.400 25.800 33.800 26.200 ;
        RECT 34.200 26.100 36.100 26.400 ;
        RECT 35.700 26.000 36.100 26.100 ;
        RECT 20.600 25.400 21.800 25.800 ;
        RECT 22.300 25.400 23.400 25.800 ;
        RECT 23.900 25.400 25.000 25.800 ;
        RECT 25.700 25.400 26.600 25.800 ;
        RECT 13.300 24.600 14.100 24.900 ;
        RECT 13.700 21.100 14.100 24.600 ;
        RECT 15.900 23.500 16.200 25.200 ;
        RECT 19.000 25.100 19.300 25.400 ;
        RECT 15.800 21.500 16.200 23.500 ;
        RECT 16.600 24.800 18.600 25.100 ;
        RECT 16.600 21.100 17.000 24.800 ;
        RECT 18.200 21.400 18.600 24.800 ;
        RECT 19.000 21.700 19.400 25.100 ;
        RECT 19.800 21.400 20.200 25.100 ;
        RECT 18.200 21.100 20.200 21.400 ;
        RECT 21.400 21.100 21.800 25.400 ;
        RECT 23.000 21.100 23.400 25.400 ;
        RECT 24.600 21.100 25.000 25.400 ;
        RECT 26.200 21.100 26.600 25.400 ;
        RECT 27.800 25.500 30.600 25.600 ;
        RECT 27.800 25.400 30.700 25.500 ;
        RECT 27.800 25.300 32.700 25.400 ;
        RECT 27.800 21.100 28.200 25.300 ;
        RECT 30.300 25.100 32.700 25.300 ;
        RECT 29.400 24.500 32.100 24.800 ;
        RECT 29.400 24.400 29.800 24.500 ;
        RECT 31.700 24.400 32.100 24.500 ;
        RECT 32.400 24.500 32.700 25.100 ;
        RECT 33.400 25.200 33.700 25.800 ;
        RECT 34.900 25.700 35.300 25.800 ;
        RECT 36.600 25.700 37.000 27.400 ;
        RECT 37.400 27.100 37.800 27.200 ;
        RECT 39.000 27.100 39.400 27.600 ;
        RECT 37.400 26.800 39.400 27.100 ;
        RECT 34.900 25.400 37.000 25.700 ;
        RECT 33.400 24.900 34.600 25.200 ;
        RECT 33.100 24.500 33.500 24.600 ;
        RECT 32.400 24.200 33.500 24.500 ;
        RECT 34.300 24.400 34.600 24.900 ;
        RECT 34.300 24.000 35.000 24.400 ;
        RECT 31.100 23.700 31.500 23.800 ;
        RECT 32.500 23.700 32.900 23.800 ;
        RECT 29.400 23.100 29.800 23.500 ;
        RECT 31.100 23.400 32.900 23.700 ;
        RECT 32.200 23.100 32.500 23.400 ;
        RECT 34.200 23.100 34.600 23.500 ;
        RECT 29.400 22.800 30.400 23.100 ;
        RECT 30.000 21.100 30.400 22.800 ;
        RECT 32.200 21.100 32.600 23.100 ;
        RECT 34.300 21.100 34.900 23.100 ;
        RECT 36.600 21.100 37.000 25.400 ;
        RECT 39.800 21.100 40.200 27.900 ;
        RECT 41.400 27.100 41.800 27.200 ;
        RECT 42.200 27.100 42.600 27.200 ;
        RECT 41.400 26.800 42.600 27.100 ;
        RECT 42.300 26.600 42.600 26.800 ;
        RECT 42.300 26.200 42.700 26.600 ;
        RECT 43.000 26.200 43.300 27.900 ;
        RECT 43.800 27.100 44.200 27.200 ;
        RECT 44.600 27.100 45.000 27.200 ;
        RECT 43.800 26.800 45.000 27.100 ;
        RECT 43.800 26.400 44.200 26.800 ;
        RECT 40.600 26.100 41.000 26.200 ;
        RECT 41.400 26.100 41.800 26.200 ;
        RECT 40.600 25.800 41.800 26.100 ;
        RECT 40.600 25.200 40.900 25.800 ;
        RECT 41.400 25.400 41.800 25.800 ;
        RECT 43.000 25.800 43.400 26.200 ;
        RECT 44.600 26.100 45.000 26.200 ;
        RECT 44.200 25.800 45.000 26.100 ;
        RECT 43.000 25.700 43.300 25.800 ;
        RECT 42.300 25.400 43.300 25.700 ;
        RECT 44.200 25.600 44.600 25.800 ;
        RECT 40.600 24.400 41.000 25.200 ;
        RECT 42.300 25.100 42.600 25.400 ;
        RECT 41.400 21.400 41.800 25.100 ;
        RECT 42.200 21.700 42.600 25.100 ;
        RECT 43.000 24.800 45.000 25.100 ;
        RECT 43.000 21.400 43.400 24.800 ;
        RECT 41.400 21.100 43.400 21.400 ;
        RECT 44.600 21.100 45.000 24.800 ;
        RECT 45.400 24.400 45.800 25.200 ;
        RECT 46.200 21.100 46.600 27.900 ;
        RECT 47.000 26.800 47.400 27.600 ;
        RECT 48.400 27.100 48.800 29.900 ;
        RECT 47.900 26.900 48.800 27.100 ;
        RECT 52.800 29.200 53.200 29.900 ;
        RECT 52.800 28.800 53.800 29.200 ;
        RECT 52.800 27.100 53.200 28.800 ;
        RECT 52.800 26.900 53.700 27.100 ;
        RECT 47.900 26.800 48.700 26.900 ;
        RECT 52.900 26.800 53.700 26.900 ;
        RECT 47.900 25.200 48.200 26.800 ;
        RECT 49.000 25.800 49.800 26.200 ;
        RECT 51.800 25.800 52.600 26.200 ;
        RECT 47.800 24.800 48.200 25.200 ;
        RECT 50.200 24.800 50.600 25.600 ;
        RECT 51.000 24.800 51.400 25.600 ;
        RECT 53.400 25.200 53.700 26.800 ;
        RECT 53.400 24.800 53.800 25.200 ;
        RECT 47.900 23.500 48.200 24.800 ;
        RECT 48.600 23.800 49.000 24.600 ;
        RECT 49.400 24.100 49.800 24.200 ;
        RECT 52.600 24.100 53.000 24.600 ;
        RECT 49.400 23.800 53.000 24.100 ;
        RECT 53.400 23.500 53.700 24.800 ;
        RECT 47.900 23.200 49.700 23.500 ;
        RECT 47.900 23.100 48.200 23.200 ;
        RECT 47.800 21.100 48.200 23.100 ;
        RECT 49.400 23.100 49.700 23.200 ;
        RECT 51.900 23.200 53.700 23.500 ;
        RECT 51.900 23.100 52.200 23.200 ;
        RECT 49.400 21.100 49.800 23.100 ;
        RECT 51.800 21.100 52.200 23.100 ;
        RECT 53.400 23.100 53.700 23.200 ;
        RECT 53.400 21.100 53.800 23.100 ;
        RECT 54.200 21.100 54.600 29.900 ;
        RECT 57.100 29.200 57.500 29.900 ;
        RECT 57.100 28.800 57.800 29.200 ;
        RECT 57.100 28.200 57.500 28.800 ;
        RECT 56.600 27.900 57.500 28.200 ;
        RECT 55.000 26.800 55.400 27.600 ;
        RECT 55.000 26.100 55.300 26.800 ;
        RECT 56.600 26.100 57.000 27.900 ;
        RECT 55.000 25.800 57.000 26.100 ;
        RECT 56.600 21.100 57.000 25.800 ;
        RECT 57.400 25.100 57.800 25.200 ;
        RECT 58.200 25.100 58.600 29.900 ;
        RECT 61.100 28.200 61.500 29.900 ;
        RECT 57.400 24.800 58.600 25.100 ;
        RECT 57.400 24.400 57.800 24.800 ;
        RECT 58.200 21.100 58.600 24.800 ;
        RECT 60.600 27.900 61.500 28.200 ;
        RECT 63.000 28.900 63.400 29.900 ;
        RECT 64.900 29.200 65.300 29.900 ;
        RECT 60.600 26.100 61.000 27.900 ;
        RECT 63.000 27.200 63.300 28.900 ;
        RECT 64.900 28.800 65.800 29.200 ;
        RECT 63.800 27.800 64.200 28.600 ;
        RECT 64.900 28.200 65.300 28.800 ;
        RECT 64.900 27.900 65.800 28.200 ;
        RECT 62.200 27.100 62.600 27.200 ;
        RECT 63.000 27.100 63.400 27.200 ;
        RECT 62.200 26.800 63.400 27.100 ;
        RECT 62.200 26.100 62.600 26.200 ;
        RECT 60.600 25.800 62.600 26.100 ;
        RECT 59.800 24.100 60.200 24.200 ;
        RECT 60.600 24.100 61.000 25.800 ;
        RECT 62.200 25.400 62.600 25.800 ;
        RECT 63.000 25.100 63.300 26.800 ;
        RECT 59.800 23.800 61.000 24.100 ;
        RECT 60.600 21.100 61.000 23.800 ;
        RECT 62.500 24.700 63.400 25.100 ;
        RECT 62.500 21.100 62.900 24.700 ;
        RECT 64.600 24.400 65.000 25.200 ;
        RECT 65.400 21.100 65.800 27.900 ;
        RECT 66.200 27.100 66.600 27.600 ;
        RECT 67.000 27.100 67.400 29.900 ;
        RECT 67.800 27.800 68.200 28.600 ;
        RECT 68.600 27.900 69.000 29.900 ;
        RECT 70.200 28.900 70.600 29.900 ;
        RECT 74.200 28.900 74.600 29.900 ;
        RECT 75.800 29.200 76.200 29.900 ;
        RECT 66.200 26.800 67.400 27.100 ;
        RECT 67.000 21.100 67.400 26.800 ;
        RECT 68.600 26.200 68.900 27.900 ;
        RECT 70.200 27.800 70.500 28.900 ;
        RECT 69.300 27.500 70.500 27.800 ;
        RECT 74.000 28.800 74.600 28.900 ;
        RECT 75.700 28.800 76.200 29.200 ;
        RECT 79.500 29.200 79.900 29.900 ;
        RECT 79.500 28.800 80.200 29.200 ;
        RECT 74.000 28.500 76.000 28.800 ;
        RECT 68.600 25.800 69.000 26.200 ;
        RECT 69.300 26.000 69.600 27.500 ;
        RECT 68.600 25.100 68.900 25.800 ;
        RECT 69.300 25.700 69.700 26.000 ;
        RECT 69.300 25.600 71.400 25.700 ;
        RECT 69.400 25.400 71.400 25.600 ;
        RECT 68.600 24.800 69.300 25.100 ;
        RECT 68.900 21.100 69.300 24.800 ;
        RECT 71.000 21.100 71.400 25.400 ;
        RECT 74.000 25.200 74.300 28.500 ;
        RECT 79.500 28.200 79.900 28.800 ;
        RECT 76.100 27.800 77.000 28.200 ;
        RECT 79.000 27.900 79.900 28.200 ;
        RECT 74.600 26.100 75.400 26.200 ;
        RECT 77.400 26.100 77.800 26.200 ;
        RECT 74.600 25.800 77.800 26.100 ;
        RECT 72.600 24.900 74.300 25.200 ;
        RECT 72.600 24.800 73.000 24.900 ;
        RECT 72.700 24.500 73.000 24.800 ;
        RECT 73.500 24.500 75.300 24.600 ;
        RECT 71.800 21.500 72.200 24.500 ;
        RECT 72.600 21.700 73.000 24.500 ;
        RECT 73.400 24.300 75.300 24.500 ;
        RECT 71.900 21.400 72.200 21.500 ;
        RECT 73.400 21.500 73.800 24.300 ;
        RECT 75.000 24.100 75.300 24.300 ;
        RECT 75.900 24.400 77.700 24.700 ;
        RECT 75.900 24.100 76.200 24.400 ;
        RECT 73.400 21.400 73.700 21.500 ;
        RECT 71.900 21.100 73.700 21.400 ;
        RECT 74.200 21.400 74.600 24.000 ;
        RECT 75.000 21.700 75.400 24.100 ;
        RECT 75.800 21.400 76.200 24.100 ;
        RECT 74.200 21.100 76.200 21.400 ;
        RECT 77.400 24.100 77.700 24.400 ;
        RECT 77.400 21.100 77.800 24.100 ;
        RECT 79.000 21.100 79.400 27.900 ;
        RECT 80.600 27.100 81.000 29.900 ;
        RECT 79.800 26.800 81.000 27.100 ;
        RECT 79.800 26.200 80.100 26.800 ;
        RECT 79.800 25.800 80.200 26.200 ;
        RECT 79.800 25.100 80.200 25.200 ;
        RECT 80.600 25.100 81.000 26.800 ;
        RECT 79.800 24.800 81.000 25.100 ;
        RECT 79.800 24.400 80.200 24.800 ;
        RECT 80.600 21.100 81.000 24.800 ;
        RECT 82.200 27.700 82.600 29.900 ;
        RECT 84.300 29.200 84.900 29.900 ;
        RECT 84.300 28.900 85.000 29.200 ;
        RECT 86.600 28.900 87.000 29.900 ;
        RECT 88.800 29.200 89.200 29.900 ;
        RECT 88.800 28.900 89.800 29.200 ;
        RECT 84.600 28.500 85.000 28.900 ;
        RECT 86.700 28.600 87.000 28.900 ;
        RECT 86.700 28.300 88.100 28.600 ;
        RECT 87.700 28.200 88.100 28.300 ;
        RECT 88.600 28.200 89.000 28.600 ;
        RECT 89.400 28.500 89.800 28.900 ;
        RECT 83.700 27.700 84.100 27.800 ;
        RECT 82.200 27.400 84.100 27.700 ;
        RECT 82.200 25.700 82.600 27.400 ;
        RECT 85.700 27.100 86.100 27.200 ;
        RECT 87.800 27.100 88.200 27.200 ;
        RECT 88.600 27.100 88.900 28.200 ;
        RECT 91.000 27.500 91.400 29.900 ;
        RECT 91.800 28.100 92.200 28.200 ;
        RECT 93.400 28.100 93.800 28.600 ;
        RECT 91.800 27.800 93.800 28.100 ;
        RECT 90.200 27.100 91.000 27.200 ;
        RECT 85.500 26.800 91.000 27.100 ;
        RECT 84.600 26.400 85.000 26.500 ;
        RECT 83.100 26.100 85.000 26.400 ;
        RECT 83.100 26.000 83.500 26.100 ;
        RECT 83.900 25.700 84.300 25.800 ;
        RECT 82.200 25.400 84.300 25.700 ;
        RECT 82.200 21.100 82.600 25.400 ;
        RECT 85.500 25.200 85.800 26.800 ;
        RECT 89.100 26.700 89.500 26.800 ;
        RECT 88.600 26.200 89.000 26.300 ;
        RECT 89.900 26.200 90.300 26.300 ;
        RECT 87.800 25.900 90.300 26.200 ;
        RECT 94.200 26.100 94.600 29.900 ;
        RECT 96.900 28.000 97.300 29.500 ;
        RECT 99.000 28.500 99.400 29.500 ;
        RECT 96.500 27.700 97.300 28.000 ;
        RECT 96.500 27.500 96.900 27.700 ;
        RECT 96.500 27.200 96.800 27.500 ;
        RECT 99.100 27.400 99.400 28.500 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 95.800 27.100 96.800 27.200 ;
        RECT 95.000 26.800 96.800 27.100 ;
        RECT 97.300 27.100 99.400 27.400 ;
        RECT 99.800 28.500 100.200 29.500 ;
        RECT 99.800 27.400 100.100 28.500 ;
        RECT 101.900 28.000 102.300 29.500 ;
        RECT 101.900 27.700 102.700 28.000 ;
        RECT 102.300 27.500 102.700 27.700 ;
        RECT 99.800 27.100 101.900 27.400 ;
        RECT 97.300 26.900 97.800 27.100 ;
        RECT 95.800 26.100 96.200 26.200 ;
        RECT 87.800 25.800 88.200 25.900 ;
        RECT 94.200 25.800 96.200 26.100 ;
        RECT 88.600 25.500 91.400 25.600 ;
        RECT 88.500 25.400 91.400 25.500 ;
        RECT 84.600 24.900 85.800 25.200 ;
        RECT 86.500 25.300 91.400 25.400 ;
        RECT 86.500 25.100 88.900 25.300 ;
        RECT 84.600 24.400 84.900 24.900 ;
        RECT 84.200 24.000 84.900 24.400 ;
        RECT 85.700 24.500 86.100 24.600 ;
        RECT 86.500 24.500 86.800 25.100 ;
        RECT 85.700 24.200 86.800 24.500 ;
        RECT 87.100 24.500 89.800 24.800 ;
        RECT 87.100 24.400 87.500 24.500 ;
        RECT 89.400 24.400 89.800 24.500 ;
        RECT 86.300 23.700 86.700 23.800 ;
        RECT 87.700 23.700 88.100 23.800 ;
        RECT 84.600 23.100 85.000 23.500 ;
        RECT 86.300 23.400 88.100 23.700 ;
        RECT 86.700 23.100 87.000 23.400 ;
        RECT 89.400 23.100 89.800 23.500 ;
        RECT 84.300 21.100 84.900 23.100 ;
        RECT 86.600 21.100 87.000 23.100 ;
        RECT 88.800 22.800 89.800 23.100 ;
        RECT 88.800 21.100 89.200 22.800 ;
        RECT 91.000 21.100 91.400 25.300 ;
        RECT 94.200 21.100 94.600 25.800 ;
        RECT 95.800 25.400 96.200 25.800 ;
        RECT 96.500 24.900 96.800 26.800 ;
        RECT 97.100 26.500 97.800 26.900 ;
        RECT 101.400 26.900 101.900 27.100 ;
        RECT 102.400 27.200 102.700 27.500 ;
        RECT 102.400 27.100 103.400 27.200 ;
        RECT 103.800 27.100 104.200 27.200 ;
        RECT 97.500 25.500 97.800 26.500 ;
        RECT 98.200 25.800 98.600 26.600 ;
        RECT 99.000 26.100 99.400 26.600 ;
        RECT 99.800 26.100 100.200 26.600 ;
        RECT 99.000 25.800 100.200 26.100 ;
        RECT 100.600 25.800 101.000 26.600 ;
        RECT 101.400 26.500 102.100 26.900 ;
        RECT 102.400 26.800 104.200 27.100 ;
        RECT 101.400 25.500 101.700 26.500 ;
        RECT 97.500 25.200 99.400 25.500 ;
        RECT 96.500 24.600 97.300 24.900 ;
        RECT 96.900 21.100 97.300 24.600 ;
        RECT 99.100 23.500 99.400 25.200 ;
        RECT 99.000 21.500 99.400 23.500 ;
        RECT 99.800 25.200 101.700 25.500 ;
        RECT 99.800 23.500 100.100 25.200 ;
        RECT 102.400 24.900 102.700 26.800 ;
        RECT 103.000 26.100 103.400 26.200 ;
        RECT 104.600 26.100 105.000 29.900 ;
        RECT 105.400 28.100 105.800 28.600 ;
        RECT 106.200 28.100 106.600 29.900 ;
        RECT 108.300 29.200 108.900 29.900 ;
        RECT 108.300 28.900 109.000 29.200 ;
        RECT 110.600 28.900 111.000 29.900 ;
        RECT 112.800 29.200 113.200 29.900 ;
        RECT 112.800 28.900 113.800 29.200 ;
        RECT 108.600 28.500 109.000 28.900 ;
        RECT 110.700 28.600 111.000 28.900 ;
        RECT 110.700 28.300 112.100 28.600 ;
        RECT 111.700 28.200 112.100 28.300 ;
        RECT 112.600 28.200 113.000 28.600 ;
        RECT 113.400 28.500 113.800 28.900 ;
        RECT 105.400 27.800 106.600 28.100 ;
        RECT 103.000 25.800 105.000 26.100 ;
        RECT 103.000 25.400 103.400 25.800 ;
        RECT 101.900 24.600 102.700 24.900 ;
        RECT 99.800 21.500 100.200 23.500 ;
        RECT 101.900 21.100 102.300 24.600 ;
        RECT 104.600 21.100 105.000 25.800 ;
        RECT 106.200 27.700 106.600 27.800 ;
        RECT 107.700 27.700 108.100 27.800 ;
        RECT 106.200 27.400 108.100 27.700 ;
        RECT 106.200 25.700 106.600 27.400 ;
        RECT 109.700 27.100 110.100 27.200 ;
        RECT 112.600 27.100 112.900 28.200 ;
        RECT 115.000 27.500 115.400 29.900 ;
        RECT 116.100 29.200 116.500 29.900 ;
        RECT 116.100 28.800 117.000 29.200 ;
        RECT 116.100 28.200 116.500 28.800 ;
        RECT 118.200 28.500 118.600 29.500 ;
        RECT 116.100 27.900 117.000 28.200 ;
        RECT 114.200 27.100 115.000 27.200 ;
        RECT 109.500 26.800 115.000 27.100 ;
        RECT 108.600 26.400 109.000 26.500 ;
        RECT 107.100 26.100 109.000 26.400 ;
        RECT 107.100 26.000 107.500 26.100 ;
        RECT 107.900 25.700 108.300 25.800 ;
        RECT 106.200 25.400 108.300 25.700 ;
        RECT 106.200 21.100 106.600 25.400 ;
        RECT 109.500 25.200 109.800 26.800 ;
        RECT 113.100 26.700 113.500 26.800 ;
        RECT 113.900 26.200 114.300 26.300 ;
        RECT 111.800 25.900 114.300 26.200 ;
        RECT 111.800 25.800 112.200 25.900 ;
        RECT 112.600 25.500 115.400 25.600 ;
        RECT 112.500 25.400 115.400 25.500 ;
        RECT 108.600 24.900 109.800 25.200 ;
        RECT 110.500 25.300 115.400 25.400 ;
        RECT 110.500 25.100 112.900 25.300 ;
        RECT 108.600 24.400 108.900 24.900 ;
        RECT 108.200 24.000 108.900 24.400 ;
        RECT 109.700 24.500 110.100 24.600 ;
        RECT 110.500 24.500 110.800 25.100 ;
        RECT 109.700 24.200 110.800 24.500 ;
        RECT 111.100 24.500 113.800 24.800 ;
        RECT 111.100 24.400 111.500 24.500 ;
        RECT 113.400 24.400 113.800 24.500 ;
        RECT 110.300 23.700 110.700 23.800 ;
        RECT 111.700 23.700 112.100 23.800 ;
        RECT 108.600 23.100 109.000 23.500 ;
        RECT 110.300 23.400 112.100 23.700 ;
        RECT 110.700 23.100 111.000 23.400 ;
        RECT 113.400 23.100 113.800 23.500 ;
        RECT 108.300 21.100 108.900 23.100 ;
        RECT 110.600 21.100 111.000 23.100 ;
        RECT 112.800 22.800 113.800 23.100 ;
        RECT 112.800 21.100 113.200 22.800 ;
        RECT 115.000 21.100 115.400 25.300 ;
        RECT 115.800 24.400 116.200 25.200 ;
        RECT 116.600 21.100 117.000 27.900 ;
        RECT 117.400 26.800 117.800 27.600 ;
        RECT 118.200 27.400 118.500 28.500 ;
        RECT 120.300 28.000 120.700 29.500 ;
        RECT 120.300 27.700 121.100 28.000 ;
        RECT 120.700 27.500 121.100 27.700 ;
        RECT 118.200 27.100 120.300 27.400 ;
        RECT 119.800 26.900 120.300 27.100 ;
        RECT 120.800 27.200 121.100 27.500 ;
        RECT 120.800 27.100 121.800 27.200 ;
        RECT 122.200 27.100 122.600 27.200 ;
        RECT 118.200 25.800 118.600 26.600 ;
        RECT 119.000 25.800 119.400 26.600 ;
        RECT 119.800 26.500 120.500 26.900 ;
        RECT 120.800 26.800 122.600 27.100 ;
        RECT 119.800 25.500 120.100 26.500 ;
        RECT 118.200 25.200 120.100 25.500 ;
        RECT 118.200 23.500 118.500 25.200 ;
        RECT 120.800 24.900 121.100 26.800 ;
        RECT 121.400 26.100 121.800 26.200 ;
        RECT 123.000 26.100 123.400 29.900 ;
        RECT 124.900 29.200 125.300 29.900 ;
        RECT 124.900 28.800 125.800 29.200 ;
        RECT 123.800 27.800 124.200 28.600 ;
        RECT 124.900 28.200 125.300 28.800 ;
        RECT 124.900 27.900 125.800 28.200 ;
        RECT 121.400 25.800 123.400 26.100 ;
        RECT 121.400 25.400 121.800 25.800 ;
        RECT 120.300 24.600 121.100 24.900 ;
        RECT 118.200 21.500 118.600 23.500 ;
        RECT 120.300 21.100 120.700 24.600 ;
        RECT 123.000 21.100 123.400 25.800 ;
        RECT 124.600 24.400 125.000 25.200 ;
        RECT 125.400 21.100 125.800 27.900 ;
        RECT 127.000 27.700 127.400 29.900 ;
        RECT 129.100 29.200 129.700 29.900 ;
        RECT 129.100 28.900 129.800 29.200 ;
        RECT 131.400 28.900 131.800 29.900 ;
        RECT 133.600 29.200 134.000 29.900 ;
        RECT 133.600 28.900 134.600 29.200 ;
        RECT 129.400 28.500 129.800 28.900 ;
        RECT 131.500 28.600 131.800 28.900 ;
        RECT 131.500 28.300 132.900 28.600 ;
        RECT 132.500 28.200 132.900 28.300 ;
        RECT 133.400 28.200 133.800 28.600 ;
        RECT 134.200 28.500 134.600 28.900 ;
        RECT 128.500 27.700 128.900 27.800 ;
        RECT 126.200 27.100 126.600 27.600 ;
        RECT 127.000 27.400 128.900 27.700 ;
        RECT 127.000 27.100 127.400 27.400 ;
        RECT 130.500 27.100 130.900 27.200 ;
        RECT 133.400 27.100 133.700 28.200 ;
        RECT 135.800 27.500 136.200 29.900 ;
        RECT 136.600 27.900 137.000 29.900 ;
        RECT 137.400 28.000 137.800 29.900 ;
        RECT 139.000 28.000 139.400 29.900 ;
        RECT 137.400 27.900 139.400 28.000 ;
        RECT 141.700 29.200 142.100 29.900 ;
        RECT 141.700 28.800 142.600 29.200 ;
        RECT 141.700 28.200 142.100 28.800 ;
        RECT 141.700 27.900 142.600 28.200 ;
        RECT 136.700 27.200 137.000 27.900 ;
        RECT 137.500 27.700 139.300 27.900 ;
        RECT 138.600 27.200 139.000 27.400 ;
        RECT 135.000 27.100 135.800 27.200 ;
        RECT 126.200 26.800 127.400 27.100 ;
        RECT 127.000 25.700 127.400 26.800 ;
        RECT 130.300 26.800 135.800 27.100 ;
        RECT 136.600 26.800 137.900 27.200 ;
        RECT 138.600 26.900 139.400 27.200 ;
        RECT 139.000 26.800 139.400 26.900 ;
        RECT 129.400 26.400 129.800 26.500 ;
        RECT 127.900 26.100 129.800 26.400 ;
        RECT 130.300 26.200 130.600 26.800 ;
        RECT 133.900 26.700 134.300 26.800 ;
        RECT 134.700 26.200 135.100 26.300 ;
        RECT 127.900 26.000 128.300 26.100 ;
        RECT 130.200 25.800 130.600 26.200 ;
        RECT 132.600 25.900 135.100 26.200 ;
        RECT 132.600 25.800 133.000 25.900 ;
        RECT 128.700 25.700 129.100 25.800 ;
        RECT 127.000 25.400 129.100 25.700 ;
        RECT 127.000 21.100 127.400 25.400 ;
        RECT 130.300 25.200 130.600 25.800 ;
        RECT 133.400 25.500 136.200 25.600 ;
        RECT 133.300 25.400 136.200 25.500 ;
        RECT 129.400 24.900 130.600 25.200 ;
        RECT 131.300 25.300 136.200 25.400 ;
        RECT 131.300 25.100 133.700 25.300 ;
        RECT 129.400 24.400 129.700 24.900 ;
        RECT 129.000 24.000 129.700 24.400 ;
        RECT 130.500 24.500 130.900 24.600 ;
        RECT 131.300 24.500 131.600 25.100 ;
        RECT 130.500 24.200 131.600 24.500 ;
        RECT 131.900 24.500 134.600 24.800 ;
        RECT 131.900 24.400 132.300 24.500 ;
        RECT 134.200 24.400 134.600 24.500 ;
        RECT 131.100 23.700 131.500 23.800 ;
        RECT 132.500 23.700 132.900 23.800 ;
        RECT 129.400 23.100 129.800 23.500 ;
        RECT 131.100 23.400 132.900 23.700 ;
        RECT 131.500 23.100 131.800 23.400 ;
        RECT 134.200 23.100 134.600 23.500 ;
        RECT 129.100 21.100 129.700 23.100 ;
        RECT 131.400 21.100 131.800 23.100 ;
        RECT 133.600 22.800 134.600 23.100 ;
        RECT 133.600 21.100 134.000 22.800 ;
        RECT 135.800 21.100 136.200 25.300 ;
        RECT 136.600 25.100 137.000 25.200 ;
        RECT 137.600 25.100 137.900 26.800 ;
        RECT 138.200 26.100 138.600 26.600 ;
        RECT 140.600 26.100 141.000 26.200 ;
        RECT 138.200 25.800 141.000 26.100 ;
        RECT 136.600 24.800 137.300 25.100 ;
        RECT 137.600 24.800 138.100 25.100 ;
        RECT 137.000 24.200 137.300 24.800 ;
        RECT 137.000 23.800 137.400 24.200 ;
        RECT 137.700 21.100 138.100 24.800 ;
        RECT 141.400 24.400 141.800 25.200 ;
        RECT 142.200 21.100 142.600 27.900 ;
        RECT 143.800 27.800 144.200 28.600 ;
        RECT 143.000 27.100 143.400 27.600 ;
        RECT 143.800 27.100 144.100 27.800 ;
        RECT 143.000 26.800 144.100 27.100 ;
        RECT 144.600 21.100 145.000 29.900 ;
        RECT 145.400 27.700 145.800 29.900 ;
        RECT 147.500 29.200 148.100 29.900 ;
        RECT 147.500 28.900 148.200 29.200 ;
        RECT 149.800 28.900 150.200 29.900 ;
        RECT 152.000 29.200 152.400 29.900 ;
        RECT 152.000 28.900 153.000 29.200 ;
        RECT 147.800 28.500 148.200 28.900 ;
        RECT 149.900 28.600 150.200 28.900 ;
        RECT 149.900 28.300 151.300 28.600 ;
        RECT 150.900 28.200 151.300 28.300 ;
        RECT 151.800 28.200 152.200 28.600 ;
        RECT 152.600 28.500 153.000 28.900 ;
        RECT 146.900 27.700 147.300 27.800 ;
        RECT 145.400 27.400 147.300 27.700 ;
        RECT 145.400 25.700 145.800 27.400 ;
        RECT 148.900 27.100 149.300 27.200 ;
        RECT 151.800 27.100 152.100 28.200 ;
        RECT 154.200 27.500 154.600 29.900 ;
        RECT 155.000 27.800 155.400 28.600 ;
        RECT 153.400 27.100 154.200 27.200 ;
        RECT 148.700 26.800 154.200 27.100 ;
        RECT 147.800 26.400 148.200 26.500 ;
        RECT 146.300 26.100 148.200 26.400 ;
        RECT 148.700 26.100 149.000 26.800 ;
        RECT 152.300 26.700 152.700 26.800 ;
        RECT 153.100 26.200 153.500 26.300 ;
        RECT 149.400 26.100 149.800 26.200 ;
        RECT 146.300 26.000 146.700 26.100 ;
        RECT 148.600 25.800 149.800 26.100 ;
        RECT 151.000 25.900 153.500 26.200 ;
        RECT 151.000 25.800 151.400 25.900 ;
        RECT 147.100 25.700 147.500 25.800 ;
        RECT 145.400 25.400 147.500 25.700 ;
        RECT 145.400 21.100 145.800 25.400 ;
        RECT 148.700 25.200 149.000 25.800 ;
        RECT 151.800 25.500 154.600 25.600 ;
        RECT 151.700 25.400 154.600 25.500 ;
        RECT 147.800 24.900 149.000 25.200 ;
        RECT 149.700 25.300 154.600 25.400 ;
        RECT 149.700 25.100 152.100 25.300 ;
        RECT 147.800 24.400 148.100 24.900 ;
        RECT 147.400 24.000 148.100 24.400 ;
        RECT 148.900 24.500 149.300 24.600 ;
        RECT 149.700 24.500 150.000 25.100 ;
        RECT 148.900 24.200 150.000 24.500 ;
        RECT 150.300 24.500 153.000 24.800 ;
        RECT 150.300 24.400 150.700 24.500 ;
        RECT 152.600 24.400 153.000 24.500 ;
        RECT 149.500 23.700 149.900 23.800 ;
        RECT 150.900 23.700 151.300 23.800 ;
        RECT 147.800 23.100 148.200 23.500 ;
        RECT 149.500 23.400 151.300 23.700 ;
        RECT 149.900 23.100 150.200 23.400 ;
        RECT 152.600 23.100 153.000 23.500 ;
        RECT 147.500 21.100 148.100 23.100 ;
        RECT 149.800 21.100 150.200 23.100 ;
        RECT 152.000 22.800 153.000 23.100 ;
        RECT 152.000 21.100 152.400 22.800 ;
        RECT 154.200 21.100 154.600 25.300 ;
        RECT 155.800 21.100 156.200 29.900 ;
        RECT 156.900 29.200 157.300 29.900 ;
        RECT 156.600 28.800 157.300 29.200 ;
        RECT 156.900 28.200 157.300 28.800 ;
        RECT 156.900 27.900 157.800 28.200 ;
        RECT 156.600 24.400 157.000 25.200 ;
        RECT 157.400 21.100 157.800 27.900 ;
        RECT 158.200 26.800 158.600 27.600 ;
        RECT 159.000 21.100 159.400 29.900 ;
        RECT 159.800 27.800 160.200 28.600 ;
        RECT 160.600 27.500 161.000 29.900 ;
        RECT 162.800 29.200 163.200 29.900 ;
        RECT 162.200 28.900 163.200 29.200 ;
        RECT 165.000 28.900 165.400 29.900 ;
        RECT 167.100 29.200 167.700 29.900 ;
        RECT 167.000 28.900 167.700 29.200 ;
        RECT 162.200 28.500 162.600 28.900 ;
        RECT 165.000 28.600 165.300 28.900 ;
        RECT 163.000 28.200 163.400 28.600 ;
        RECT 163.900 28.300 165.300 28.600 ;
        RECT 167.000 28.500 167.400 28.900 ;
        RECT 163.900 28.200 164.300 28.300 ;
        RECT 161.000 27.100 161.800 27.200 ;
        RECT 163.100 27.100 163.400 28.200 ;
        RECT 167.900 27.700 168.300 27.800 ;
        RECT 169.400 27.700 169.800 29.900 ;
        RECT 167.900 27.400 169.800 27.700 ;
        RECT 165.900 27.100 166.300 27.200 ;
        RECT 161.000 26.800 166.500 27.100 ;
        RECT 162.500 26.700 162.900 26.800 ;
        RECT 161.700 26.200 162.100 26.300 ;
        RECT 161.700 26.100 164.200 26.200 ;
        RECT 164.600 26.100 165.000 26.200 ;
        RECT 161.700 25.900 165.000 26.100 ;
        RECT 163.800 25.800 165.000 25.900 ;
        RECT 160.600 25.500 163.400 25.600 ;
        RECT 160.600 25.400 163.500 25.500 ;
        RECT 160.600 25.300 165.500 25.400 ;
        RECT 160.600 21.100 161.000 25.300 ;
        RECT 163.100 25.100 165.500 25.300 ;
        RECT 162.200 24.500 164.900 24.800 ;
        RECT 162.200 24.400 162.600 24.500 ;
        RECT 164.500 24.400 164.900 24.500 ;
        RECT 165.200 24.500 165.500 25.100 ;
        RECT 166.200 25.200 166.500 26.800 ;
        RECT 167.000 26.400 167.400 26.500 ;
        RECT 167.000 26.100 168.900 26.400 ;
        RECT 168.500 26.000 168.900 26.100 ;
        RECT 167.700 25.700 168.100 25.800 ;
        RECT 169.400 25.700 169.800 27.400 ;
        RECT 167.700 25.400 169.800 25.700 ;
        RECT 166.200 24.900 167.400 25.200 ;
        RECT 165.900 24.500 166.300 24.600 ;
        RECT 165.200 24.200 166.300 24.500 ;
        RECT 167.100 24.400 167.400 24.900 ;
        RECT 167.100 24.000 167.800 24.400 ;
        RECT 163.900 23.700 164.300 23.800 ;
        RECT 165.300 23.700 165.700 23.800 ;
        RECT 162.200 23.100 162.600 23.500 ;
        RECT 163.900 23.400 165.700 23.700 ;
        RECT 165.000 23.100 165.300 23.400 ;
        RECT 167.000 23.100 167.400 23.500 ;
        RECT 162.200 22.800 163.200 23.100 ;
        RECT 162.800 21.100 163.200 22.800 ;
        RECT 165.000 21.100 165.400 23.100 ;
        RECT 167.100 21.100 167.700 23.100 ;
        RECT 169.400 21.100 169.800 25.400 ;
        RECT 170.200 21.100 170.600 29.900 ;
        RECT 171.000 27.800 171.400 28.600 ;
        RECT 171.800 27.900 172.200 29.900 ;
        RECT 172.600 28.000 173.000 29.900 ;
        RECT 174.200 28.000 174.600 29.900 ;
        RECT 172.600 27.900 174.600 28.000 ;
        RECT 175.000 28.000 175.400 29.900 ;
        RECT 176.600 28.000 177.000 29.900 ;
        RECT 175.000 27.900 177.000 28.000 ;
        RECT 177.400 27.900 177.800 29.900 ;
        RECT 178.500 28.200 178.900 29.900 ;
        RECT 178.500 27.900 179.400 28.200 ;
        RECT 171.900 27.200 172.200 27.900 ;
        RECT 172.700 27.700 174.500 27.900 ;
        RECT 175.100 27.700 176.900 27.900 ;
        RECT 173.800 27.200 174.200 27.400 ;
        RECT 175.400 27.200 175.800 27.400 ;
        RECT 177.400 27.200 177.700 27.900 ;
        RECT 171.800 26.800 173.100 27.200 ;
        RECT 173.800 27.100 174.600 27.200 ;
        RECT 175.000 27.100 175.800 27.200 ;
        RECT 173.800 26.900 175.800 27.100 ;
        RECT 174.200 26.800 175.400 26.900 ;
        RECT 176.500 26.800 177.800 27.200 ;
        RECT 171.800 25.100 172.200 25.200 ;
        RECT 172.800 25.100 173.100 26.800 ;
        RECT 173.400 25.800 173.800 26.600 ;
        RECT 175.800 25.800 176.200 26.600 ;
        RECT 176.500 25.100 176.800 26.800 ;
        RECT 179.000 26.100 179.400 27.900 ;
        RECT 179.800 26.800 180.200 27.600 ;
        RECT 177.400 25.800 179.400 26.100 ;
        RECT 177.400 25.200 177.700 25.800 ;
        RECT 177.400 25.100 177.800 25.200 ;
        RECT 171.800 24.800 172.500 25.100 ;
        RECT 172.800 24.800 173.300 25.100 ;
        RECT 172.200 24.200 172.500 24.800 ;
        RECT 172.200 23.800 172.600 24.200 ;
        RECT 172.900 21.100 173.300 24.800 ;
        RECT 176.300 24.800 176.800 25.100 ;
        RECT 177.100 24.800 177.800 25.100 ;
        RECT 176.300 21.100 176.700 24.800 ;
        RECT 177.100 24.200 177.400 24.800 ;
        RECT 178.200 24.400 178.600 25.200 ;
        RECT 177.000 23.800 177.400 24.200 ;
        RECT 179.000 21.100 179.400 25.800 ;
        RECT 2.500 16.400 2.900 19.900 ;
        RECT 4.600 17.500 5.000 19.500 ;
        RECT 2.100 16.100 2.900 16.400 ;
        RECT 1.400 14.800 1.800 15.600 ;
        RECT 2.100 14.200 2.400 16.100 ;
        RECT 4.700 15.800 5.000 17.500 ;
        RECT 3.100 15.500 5.000 15.800 ;
        RECT 5.400 16.100 5.800 19.900 ;
        RECT 7.000 16.200 7.400 19.900 ;
        RECT 8.600 16.200 9.000 19.900 ;
        RECT 6.200 16.100 6.600 16.200 ;
        RECT 5.400 15.800 6.600 16.100 ;
        RECT 7.000 15.900 9.000 16.200 ;
        RECT 9.400 15.900 9.800 19.900 ;
        RECT 10.500 16.300 10.900 19.900 ;
        RECT 10.500 15.900 11.400 16.300 ;
        RECT 3.100 14.500 3.400 15.500 ;
        RECT 1.400 13.800 2.400 14.200 ;
        RECT 2.700 14.100 3.400 14.500 ;
        RECT 3.800 14.400 4.200 15.200 ;
        RECT 4.600 14.400 5.000 15.200 ;
        RECT 2.100 13.500 2.400 13.800 ;
        RECT 2.900 13.900 3.400 14.100 ;
        RECT 2.900 13.600 5.000 13.900 ;
        RECT 2.100 13.300 2.500 13.500 ;
        RECT 2.100 13.000 2.900 13.300 ;
        RECT 2.500 12.200 2.900 13.000 ;
        RECT 4.700 12.500 5.000 13.600 ;
        RECT 2.500 11.800 3.400 12.200 ;
        RECT 2.500 11.500 2.900 11.800 ;
        RECT 4.600 11.500 5.000 12.500 ;
        RECT 5.400 11.100 5.800 15.800 ;
        RECT 7.400 15.200 7.800 15.400 ;
        RECT 9.400 15.200 9.700 15.900 ;
        RECT 7.000 14.900 7.800 15.200 ;
        RECT 8.600 14.900 9.800 15.200 ;
        RECT 7.000 14.800 7.400 14.900 ;
        RECT 7.800 13.800 8.200 14.600 ;
        RECT 6.200 12.400 6.600 13.200 ;
        RECT 8.600 13.100 8.900 14.900 ;
        RECT 9.400 14.800 9.800 14.900 ;
        RECT 10.200 14.800 10.600 15.600 ;
        RECT 11.000 14.200 11.300 15.900 ;
        RECT 12.600 15.600 13.000 19.900 ;
        RECT 14.700 17.900 15.300 19.900 ;
        RECT 17.000 17.900 17.400 19.900 ;
        RECT 19.200 18.200 19.600 19.900 ;
        RECT 19.200 17.900 20.200 18.200 ;
        RECT 15.000 17.500 15.400 17.900 ;
        RECT 17.100 17.600 17.400 17.900 ;
        RECT 16.700 17.300 18.500 17.600 ;
        RECT 19.800 17.500 20.200 17.900 ;
        RECT 16.700 17.200 17.100 17.300 ;
        RECT 18.100 17.200 18.500 17.300 ;
        RECT 14.200 17.000 14.900 17.200 ;
        RECT 14.200 16.800 15.300 17.000 ;
        RECT 14.600 16.600 15.300 16.800 ;
        RECT 15.000 16.100 15.300 16.600 ;
        RECT 16.100 16.500 17.200 16.800 ;
        RECT 16.100 16.400 16.500 16.500 ;
        RECT 15.000 15.800 16.200 16.100 ;
        RECT 12.600 15.300 14.700 15.600 ;
        RECT 11.000 13.800 11.400 14.200 ;
        RECT 9.400 13.100 9.800 13.200 ;
        RECT 11.000 13.100 11.300 13.800 ;
        RECT 12.600 13.600 13.000 15.300 ;
        RECT 14.300 15.200 14.700 15.300 ;
        RECT 13.500 14.900 13.900 15.000 ;
        RECT 13.500 14.600 15.400 14.900 ;
        RECT 15.000 14.500 15.400 14.600 ;
        RECT 15.900 14.200 16.200 15.800 ;
        RECT 16.900 15.900 17.200 16.500 ;
        RECT 17.500 16.500 17.900 16.600 ;
        RECT 19.800 16.500 20.200 16.600 ;
        RECT 17.500 16.200 20.200 16.500 ;
        RECT 16.900 15.700 19.300 15.900 ;
        RECT 21.400 15.700 21.800 19.900 ;
        RECT 16.900 15.600 21.800 15.700 ;
        RECT 18.900 15.500 21.800 15.600 ;
        RECT 22.200 17.500 22.600 19.500 ;
        RECT 22.200 15.800 22.500 17.500 ;
        RECT 24.300 16.400 24.700 19.900 ;
        RECT 24.300 16.100 25.100 16.400 ;
        RECT 22.200 15.500 24.100 15.800 ;
        RECT 19.000 15.400 21.800 15.500 ;
        RECT 18.200 15.100 18.600 15.200 ;
        RECT 18.200 14.800 20.700 15.100 ;
        RECT 19.000 14.700 19.400 14.800 ;
        RECT 20.300 14.700 20.700 14.800 ;
        RECT 22.200 14.400 22.600 15.200 ;
        RECT 23.000 14.400 23.400 15.200 ;
        RECT 23.800 14.500 24.100 15.500 ;
        RECT 19.500 14.200 19.900 14.300 ;
        RECT 15.900 13.900 21.400 14.200 ;
        RECT 23.800 14.100 24.500 14.500 ;
        RECT 24.800 14.200 25.100 16.100 ;
        RECT 25.400 15.100 25.800 15.600 ;
        RECT 27.000 15.100 27.400 19.900 ;
        RECT 28.600 15.700 29.000 19.900 ;
        RECT 30.800 18.200 31.200 19.900 ;
        RECT 30.200 17.900 31.200 18.200 ;
        RECT 33.000 17.900 33.400 19.900 ;
        RECT 35.100 17.900 35.700 19.900 ;
        RECT 30.200 17.500 30.600 17.900 ;
        RECT 33.000 17.600 33.300 17.900 ;
        RECT 31.900 17.300 33.700 17.600 ;
        RECT 35.000 17.500 35.400 17.900 ;
        RECT 31.900 17.200 32.300 17.300 ;
        RECT 33.300 17.200 33.700 17.300 ;
        RECT 30.200 16.500 30.600 16.600 ;
        RECT 32.500 16.500 32.900 16.600 ;
        RECT 30.200 16.200 32.900 16.500 ;
        RECT 33.200 16.500 34.300 16.800 ;
        RECT 33.200 15.900 33.500 16.500 ;
        RECT 33.900 16.400 34.300 16.500 ;
        RECT 35.100 16.600 35.800 17.000 ;
        RECT 35.100 16.100 35.400 16.600 ;
        RECT 31.100 15.700 33.500 15.900 ;
        RECT 28.600 15.600 33.500 15.700 ;
        RECT 34.200 15.800 35.400 16.100 ;
        RECT 28.600 15.500 31.500 15.600 ;
        RECT 28.600 15.400 31.400 15.500 ;
        RECT 31.800 15.100 32.200 15.200 ;
        RECT 25.400 14.800 27.400 15.100 ;
        RECT 23.800 13.900 24.300 14.100 ;
        RECT 16.100 13.800 16.500 13.900 ;
        RECT 18.200 13.800 18.600 13.900 ;
        RECT 12.600 13.300 14.600 13.600 ;
        RECT 8.600 11.100 9.000 13.100 ;
        RECT 9.400 12.800 11.300 13.100 ;
        RECT 9.300 12.400 9.700 12.800 ;
        RECT 11.000 12.100 11.300 12.800 ;
        RECT 11.800 12.400 12.200 13.200 ;
        RECT 11.000 11.100 11.400 12.100 ;
        RECT 12.600 11.100 13.000 13.300 ;
        RECT 14.100 13.200 14.600 13.300 ;
        RECT 14.200 13.100 14.600 13.200 ;
        RECT 15.800 13.100 16.200 13.200 ;
        RECT 14.200 12.800 16.200 13.100 ;
        RECT 19.000 12.800 19.300 13.900 ;
        RECT 20.600 13.800 21.400 13.900 ;
        RECT 22.200 13.600 24.300 13.900 ;
        RECT 24.800 13.800 25.800 14.200 ;
        RECT 18.100 12.700 18.500 12.800 ;
        RECT 15.000 12.100 15.400 12.500 ;
        RECT 17.100 12.400 18.500 12.700 ;
        RECT 19.000 12.400 19.400 12.800 ;
        RECT 17.100 12.100 17.400 12.400 ;
        RECT 19.800 12.100 20.200 12.500 ;
        RECT 14.700 11.800 15.400 12.100 ;
        RECT 14.700 11.100 15.300 11.800 ;
        RECT 17.000 11.100 17.400 12.100 ;
        RECT 19.200 11.800 20.200 12.100 ;
        RECT 19.200 11.100 19.600 11.800 ;
        RECT 21.400 11.100 21.800 13.500 ;
        RECT 22.200 12.500 22.500 13.600 ;
        RECT 24.800 13.500 25.100 13.800 ;
        RECT 24.700 13.300 25.100 13.500 ;
        RECT 24.300 13.000 25.100 13.300 ;
        RECT 22.200 11.500 22.600 12.500 ;
        RECT 24.300 12.200 24.700 13.000 ;
        RECT 24.300 11.800 25.000 12.200 ;
        RECT 24.300 11.500 24.700 11.800 ;
        RECT 27.000 11.100 27.400 14.800 ;
        RECT 29.700 14.800 32.200 15.100 ;
        RECT 33.400 15.100 33.800 15.200 ;
        RECT 34.200 15.100 34.500 15.800 ;
        RECT 37.400 15.600 37.800 19.900 ;
        RECT 35.700 15.300 37.800 15.600 ;
        RECT 39.800 17.500 40.200 19.500 ;
        RECT 39.800 15.800 40.100 17.500 ;
        RECT 41.900 16.400 42.300 19.900 ;
        RECT 41.900 16.100 42.700 16.400 ;
        RECT 39.800 15.500 41.700 15.800 ;
        RECT 35.700 15.200 36.100 15.300 ;
        RECT 33.400 14.800 34.500 15.100 ;
        RECT 36.500 14.900 36.900 15.000 ;
        RECT 29.700 14.700 30.100 14.800 ;
        RECT 30.500 14.200 30.900 14.300 ;
        RECT 34.200 14.200 34.500 14.800 ;
        RECT 35.000 14.600 36.900 14.900 ;
        RECT 35.000 14.500 35.400 14.600 ;
        RECT 29.000 13.900 34.500 14.200 ;
        RECT 29.000 13.800 29.800 13.900 ;
        RECT 27.800 12.400 28.200 13.200 ;
        RECT 28.600 11.100 29.000 13.500 ;
        RECT 31.100 12.800 31.400 13.900 ;
        RECT 33.900 13.800 34.300 13.900 ;
        RECT 37.400 13.600 37.800 15.300 ;
        RECT 39.800 14.400 40.200 15.200 ;
        RECT 40.600 14.400 41.000 15.200 ;
        RECT 41.400 14.500 41.700 15.500 ;
        RECT 41.400 14.100 42.100 14.500 ;
        RECT 42.400 14.200 42.700 16.100 ;
        RECT 43.000 15.100 43.400 15.600 ;
        RECT 45.400 15.100 45.800 19.900 ;
        RECT 43.000 14.800 45.800 15.100 ;
        RECT 41.400 13.900 41.900 14.100 ;
        RECT 35.900 13.300 37.800 13.600 ;
        RECT 35.900 13.200 36.300 13.300 ;
        RECT 30.200 12.100 30.600 12.500 ;
        RECT 31.000 12.400 31.400 12.800 ;
        RECT 31.900 12.700 32.300 12.800 ;
        RECT 31.900 12.400 33.300 12.700 ;
        RECT 33.000 12.100 33.300 12.400 ;
        RECT 35.000 12.100 35.400 12.500 ;
        RECT 30.200 11.800 31.200 12.100 ;
        RECT 30.800 11.100 31.200 11.800 ;
        RECT 33.000 11.100 33.400 12.100 ;
        RECT 35.000 11.800 35.700 12.100 ;
        RECT 35.100 11.100 35.700 11.800 ;
        RECT 37.400 11.100 37.800 13.300 ;
        RECT 39.800 13.600 41.900 13.900 ;
        RECT 42.400 13.800 43.400 14.200 ;
        RECT 44.600 13.800 45.000 14.200 ;
        RECT 39.800 12.500 40.100 13.600 ;
        RECT 42.400 13.500 42.700 13.800 ;
        RECT 42.300 13.300 42.700 13.500 ;
        RECT 41.900 13.200 42.700 13.300 ;
        RECT 41.400 13.000 42.700 13.200 ;
        RECT 44.600 13.200 44.900 13.800 ;
        RECT 41.400 12.800 42.300 13.000 ;
        RECT 39.800 11.500 40.200 12.500 ;
        RECT 41.900 11.500 42.300 12.800 ;
        RECT 44.600 12.400 45.000 13.200 ;
        RECT 45.400 11.100 45.800 14.800 ;
        RECT 46.200 15.600 46.600 19.900 ;
        RECT 48.300 17.900 48.900 19.900 ;
        RECT 50.600 17.900 51.000 19.900 ;
        RECT 52.800 18.200 53.200 19.900 ;
        RECT 52.800 17.900 53.800 18.200 ;
        RECT 48.600 17.500 49.000 17.900 ;
        RECT 50.700 17.600 51.000 17.900 ;
        RECT 50.300 17.300 52.100 17.600 ;
        RECT 53.400 17.500 53.800 17.900 ;
        RECT 50.300 17.200 50.700 17.300 ;
        RECT 51.700 17.200 52.100 17.300 ;
        RECT 48.200 16.600 48.900 17.000 ;
        RECT 48.600 16.100 48.900 16.600 ;
        RECT 49.700 16.500 50.800 16.800 ;
        RECT 49.700 16.400 50.100 16.500 ;
        RECT 48.600 15.800 49.800 16.100 ;
        RECT 46.200 15.300 48.300 15.600 ;
        RECT 46.200 13.600 46.600 15.300 ;
        RECT 47.900 15.200 48.300 15.300 ;
        RECT 47.100 14.900 47.500 15.000 ;
        RECT 47.100 14.600 49.000 14.900 ;
        RECT 48.600 14.500 49.000 14.600 ;
        RECT 49.500 14.200 49.800 15.800 ;
        RECT 50.500 15.900 50.800 16.500 ;
        RECT 51.100 16.500 51.500 16.600 ;
        RECT 53.400 16.500 53.800 16.600 ;
        RECT 51.100 16.200 53.800 16.500 ;
        RECT 50.500 15.700 52.900 15.900 ;
        RECT 55.000 15.700 55.400 19.900 ;
        RECT 57.100 16.300 57.500 19.900 ;
        RECT 56.600 15.900 57.500 16.300 ;
        RECT 58.200 15.900 58.600 19.900 ;
        RECT 59.000 16.200 59.400 19.900 ;
        RECT 60.600 16.200 61.000 19.900 ;
        RECT 59.000 15.900 61.000 16.200 ;
        RECT 50.500 15.600 55.400 15.700 ;
        RECT 52.500 15.500 55.400 15.600 ;
        RECT 52.600 15.400 55.400 15.500 ;
        RECT 51.800 15.100 52.200 15.200 ;
        RECT 51.800 14.800 54.300 15.100 ;
        RECT 52.600 14.700 53.000 14.800 ;
        RECT 53.900 14.700 54.300 14.800 ;
        RECT 53.100 14.200 53.500 14.300 ;
        RECT 56.700 14.200 57.000 15.900 ;
        RECT 57.400 14.800 57.800 15.600 ;
        RECT 58.300 15.200 58.600 15.900 ;
        RECT 60.200 15.200 60.600 15.400 ;
        RECT 58.200 14.900 59.400 15.200 ;
        RECT 60.200 14.900 61.000 15.200 ;
        RECT 58.200 14.800 58.600 14.900 ;
        RECT 49.500 13.900 55.000 14.200 ;
        RECT 49.700 13.800 50.100 13.900 ;
        RECT 46.200 13.300 48.200 13.600 ;
        RECT 46.200 11.100 46.600 13.300 ;
        RECT 47.700 13.200 48.200 13.300 ;
        RECT 52.600 13.200 52.900 13.900 ;
        RECT 54.200 13.800 55.000 13.900 ;
        RECT 56.600 13.800 57.000 14.200 ;
        RECT 47.800 13.100 48.200 13.200 ;
        RECT 49.400 13.100 49.800 13.200 ;
        RECT 47.800 12.800 49.800 13.100 ;
        RECT 51.700 12.700 52.100 12.800 ;
        RECT 48.600 12.100 49.000 12.500 ;
        RECT 50.700 12.400 52.100 12.700 ;
        RECT 52.600 12.400 53.000 13.200 ;
        RECT 50.700 12.100 51.000 12.400 ;
        RECT 53.400 12.100 53.800 12.500 ;
        RECT 48.300 11.800 49.000 12.100 ;
        RECT 48.300 11.100 48.900 11.800 ;
        RECT 50.600 11.100 51.000 12.100 ;
        RECT 52.800 11.800 53.800 12.100 ;
        RECT 52.800 11.100 53.200 11.800 ;
        RECT 55.000 11.100 55.400 13.500 ;
        RECT 55.800 12.400 56.200 13.200 ;
        RECT 56.700 13.100 57.000 13.800 ;
        RECT 59.100 13.200 59.400 14.900 ;
        RECT 60.600 14.800 61.000 14.900 ;
        RECT 62.200 15.100 62.600 19.900 ;
        RECT 64.900 16.400 65.300 19.900 ;
        RECT 67.000 17.500 67.400 19.500 ;
        RECT 64.500 16.100 65.300 16.400 ;
        RECT 63.800 15.100 64.200 15.600 ;
        RECT 62.200 14.800 64.200 15.100 ;
        RECT 59.800 13.800 60.200 14.600 ;
        RECT 58.200 13.100 58.600 13.200 ;
        RECT 56.600 12.800 58.600 13.100 ;
        RECT 56.700 12.100 57.000 12.800 ;
        RECT 58.300 12.400 58.700 12.800 ;
        RECT 56.600 11.100 57.000 12.100 ;
        RECT 59.000 11.100 59.400 13.200 ;
        RECT 61.400 12.400 61.800 13.200 ;
        RECT 62.200 11.100 62.600 14.800 ;
        RECT 64.500 14.200 64.800 16.100 ;
        RECT 67.100 15.800 67.400 17.500 ;
        RECT 67.800 15.800 68.200 16.600 ;
        RECT 65.500 15.500 67.400 15.800 ;
        RECT 65.500 14.500 65.800 15.500 ;
        RECT 63.000 14.100 63.400 14.200 ;
        RECT 63.800 14.100 64.800 14.200 ;
        RECT 65.100 14.100 65.800 14.500 ;
        RECT 66.200 14.400 66.600 15.200 ;
        RECT 67.000 14.400 67.400 15.200 ;
        RECT 63.000 13.800 64.800 14.100 ;
        RECT 64.500 13.500 64.800 13.800 ;
        RECT 65.300 13.900 65.800 14.100 ;
        RECT 65.300 13.600 67.400 13.900 ;
        RECT 64.500 13.300 64.900 13.500 ;
        RECT 64.500 13.000 65.300 13.300 ;
        RECT 64.900 11.500 65.300 13.000 ;
        RECT 67.100 12.500 67.400 13.600 ;
        RECT 68.600 13.100 69.000 19.900 ;
        RECT 71.500 16.300 71.900 19.900 ;
        RECT 71.000 15.900 71.900 16.300 ;
        RECT 72.600 15.900 73.000 19.900 ;
        RECT 73.400 16.200 73.800 19.900 ;
        RECT 75.000 16.200 75.400 19.900 ;
        RECT 73.400 15.900 75.400 16.200 ;
        RECT 71.100 14.200 71.400 15.900 ;
        RECT 71.800 14.800 72.200 15.600 ;
        RECT 72.700 15.200 73.000 15.900 ;
        RECT 76.600 15.600 77.000 19.900 ;
        RECT 78.200 15.600 78.600 19.900 ;
        RECT 74.600 15.200 75.000 15.400 ;
        RECT 76.600 15.200 78.600 15.600 ;
        RECT 79.800 15.600 80.200 19.900 ;
        RECT 81.900 17.900 82.500 19.900 ;
        RECT 84.200 17.900 84.600 19.900 ;
        RECT 86.400 18.200 86.800 19.900 ;
        RECT 86.400 17.900 87.400 18.200 ;
        RECT 82.200 17.500 82.600 17.900 ;
        RECT 84.300 17.600 84.600 17.900 ;
        RECT 83.900 17.300 85.700 17.600 ;
        RECT 87.000 17.500 87.400 17.900 ;
        RECT 83.900 17.200 84.300 17.300 ;
        RECT 85.300 17.200 85.700 17.300 ;
        RECT 81.800 16.600 82.500 17.000 ;
        RECT 82.200 16.100 82.500 16.600 ;
        RECT 83.300 16.500 84.400 16.800 ;
        RECT 83.300 16.400 83.700 16.500 ;
        RECT 82.200 15.800 83.400 16.100 ;
        RECT 79.800 15.300 81.900 15.600 ;
        RECT 72.600 14.900 73.800 15.200 ;
        RECT 74.600 14.900 75.400 15.200 ;
        RECT 72.600 14.800 73.000 14.900 ;
        RECT 69.400 14.100 69.800 14.200 ;
        RECT 69.400 13.800 70.500 14.100 ;
        RECT 71.000 13.800 71.400 14.200 ;
        RECT 69.400 13.400 69.800 13.800 ;
        RECT 67.000 11.500 67.400 12.500 ;
        RECT 68.100 12.800 69.000 13.100 ;
        RECT 70.200 13.200 70.500 13.800 ;
        RECT 68.100 11.100 68.500 12.800 ;
        RECT 70.200 12.400 70.600 13.200 ;
        RECT 71.100 13.100 71.400 13.800 ;
        RECT 72.600 13.100 73.000 13.200 ;
        RECT 73.500 13.100 73.800 14.900 ;
        RECT 75.000 14.800 75.400 14.900 ;
        RECT 74.200 13.800 74.600 14.600 ;
        RECT 76.600 13.800 77.000 15.200 ;
        RECT 71.000 12.800 73.000 13.100 ;
        RECT 71.100 12.100 71.400 12.800 ;
        RECT 72.700 12.400 73.100 12.800 ;
        RECT 71.000 11.100 71.400 12.100 ;
        RECT 73.400 11.100 73.800 13.100 ;
        RECT 76.600 13.400 78.600 13.800 ;
        RECT 76.600 11.100 77.000 13.400 ;
        RECT 78.200 11.100 78.600 13.400 ;
        RECT 79.800 13.600 80.200 15.300 ;
        RECT 81.500 15.200 81.900 15.300 ;
        RECT 80.700 14.900 81.100 15.000 ;
        RECT 80.700 14.600 82.600 14.900 ;
        RECT 82.200 14.500 82.600 14.600 ;
        RECT 83.100 14.200 83.400 15.800 ;
        RECT 84.100 15.900 84.400 16.500 ;
        RECT 84.700 16.500 85.100 16.600 ;
        RECT 87.000 16.500 87.400 16.600 ;
        RECT 84.700 16.200 87.400 16.500 ;
        RECT 84.100 15.700 86.500 15.900 ;
        RECT 88.600 15.700 89.000 19.900 ;
        RECT 84.100 15.600 89.000 15.700 ;
        RECT 86.100 15.500 89.000 15.600 ;
        RECT 86.200 15.400 89.000 15.500 ;
        RECT 85.400 15.100 85.800 15.200 ;
        RECT 91.800 15.100 92.200 19.900 ;
        RECT 94.500 16.400 94.900 19.900 ;
        RECT 96.600 17.500 97.000 19.500 ;
        RECT 94.100 16.100 94.900 16.400 ;
        RECT 93.400 15.100 93.800 15.600 ;
        RECT 85.400 14.800 87.900 15.100 ;
        RECT 86.200 14.700 86.600 14.800 ;
        RECT 87.500 14.700 87.900 14.800 ;
        RECT 91.800 14.800 93.800 15.100 ;
        RECT 86.700 14.200 87.100 14.300 ;
        RECT 83.000 13.900 88.600 14.200 ;
        RECT 83.000 13.800 83.700 13.900 ;
        RECT 79.800 13.300 81.700 13.600 ;
        RECT 79.800 11.100 80.200 13.300 ;
        RECT 81.300 13.200 81.700 13.300 ;
        RECT 86.200 12.800 86.500 13.900 ;
        RECT 87.800 13.800 88.600 13.900 ;
        RECT 85.300 12.700 85.700 12.800 ;
        RECT 82.200 12.100 82.600 12.500 ;
        RECT 84.300 12.400 85.700 12.700 ;
        RECT 86.200 12.400 86.600 12.800 ;
        RECT 84.300 12.100 84.600 12.400 ;
        RECT 87.000 12.100 87.400 12.500 ;
        RECT 81.900 11.800 82.600 12.100 ;
        RECT 81.900 11.100 82.500 11.800 ;
        RECT 84.200 11.100 84.600 12.100 ;
        RECT 86.400 11.800 87.400 12.100 ;
        RECT 86.400 11.100 86.800 11.800 ;
        RECT 88.600 11.100 89.000 13.500 ;
        RECT 91.000 12.400 91.400 13.200 ;
        RECT 91.800 11.100 92.200 14.800 ;
        RECT 94.100 14.200 94.400 16.100 ;
        RECT 96.700 15.800 97.000 17.500 ;
        RECT 95.100 15.500 97.000 15.800 ;
        RECT 97.400 15.600 97.800 19.900 ;
        RECT 99.500 17.900 100.100 19.900 ;
        RECT 101.800 17.900 102.200 19.900 ;
        RECT 104.000 18.200 104.400 19.900 ;
        RECT 104.000 17.900 105.000 18.200 ;
        RECT 99.800 17.500 100.200 17.900 ;
        RECT 101.900 17.600 102.200 17.900 ;
        RECT 101.500 17.300 103.300 17.600 ;
        RECT 104.600 17.500 105.000 17.900 ;
        RECT 101.500 17.200 101.900 17.300 ;
        RECT 102.900 17.200 103.300 17.300 ;
        RECT 99.400 16.600 100.100 17.000 ;
        RECT 99.800 16.100 100.100 16.600 ;
        RECT 100.900 16.500 102.000 16.800 ;
        RECT 100.900 16.400 101.300 16.500 ;
        RECT 99.800 15.800 101.000 16.100 ;
        RECT 95.100 14.500 95.400 15.500 ;
        RECT 97.400 15.300 99.500 15.600 ;
        RECT 92.600 14.100 93.000 14.200 ;
        RECT 93.400 14.100 94.400 14.200 ;
        RECT 94.700 14.100 95.400 14.500 ;
        RECT 95.800 14.400 96.200 15.200 ;
        RECT 96.600 14.400 97.000 15.200 ;
        RECT 92.600 13.800 94.400 14.100 ;
        RECT 94.100 13.500 94.400 13.800 ;
        RECT 94.900 13.900 95.400 14.100 ;
        RECT 94.900 13.600 97.000 13.900 ;
        RECT 94.100 13.300 94.500 13.500 ;
        RECT 94.100 13.000 94.900 13.300 ;
        RECT 94.500 11.500 94.900 13.000 ;
        RECT 96.700 12.500 97.000 13.600 ;
        RECT 96.600 11.500 97.000 12.500 ;
        RECT 97.400 13.600 97.800 15.300 ;
        RECT 99.100 15.200 99.500 15.300 ;
        RECT 100.700 15.200 101.000 15.800 ;
        RECT 101.700 15.900 102.000 16.500 ;
        RECT 102.300 16.500 102.700 16.600 ;
        RECT 104.600 16.500 105.000 16.600 ;
        RECT 102.300 16.200 105.000 16.500 ;
        RECT 101.700 15.700 104.100 15.900 ;
        RECT 106.200 15.700 106.600 19.900 ;
        RECT 101.700 15.600 106.600 15.700 ;
        RECT 103.700 15.500 106.600 15.600 ;
        RECT 103.800 15.400 106.600 15.500 ;
        RECT 98.300 14.900 98.700 15.000 ;
        RECT 98.300 14.600 100.200 14.900 ;
        RECT 100.600 14.800 101.000 15.200 ;
        RECT 103.000 15.100 103.400 15.200 ;
        RECT 107.800 15.100 108.200 19.900 ;
        RECT 110.500 16.400 110.900 19.900 ;
        RECT 112.600 17.500 113.000 19.500 ;
        RECT 110.100 16.100 110.900 16.400 ;
        RECT 110.100 15.800 110.600 16.100 ;
        RECT 112.700 15.800 113.000 17.500 ;
        RECT 113.400 16.100 113.800 16.200 ;
        RECT 114.200 16.100 114.600 19.900 ;
        RECT 113.400 15.800 114.600 16.100 ;
        RECT 109.400 15.100 109.800 15.600 ;
        RECT 103.000 14.800 105.500 15.100 ;
        RECT 99.800 14.500 100.200 14.600 ;
        RECT 100.700 14.200 101.000 14.800 ;
        RECT 103.800 14.700 104.200 14.800 ;
        RECT 105.100 14.700 105.500 14.800 ;
        RECT 107.800 14.800 109.800 15.100 ;
        RECT 104.300 14.200 104.700 14.300 ;
        RECT 100.700 13.900 106.200 14.200 ;
        RECT 100.900 13.800 101.300 13.900 ;
        RECT 97.400 13.300 99.300 13.600 ;
        RECT 97.400 11.100 97.800 13.300 ;
        RECT 98.900 13.200 99.300 13.300 ;
        RECT 103.800 12.800 104.100 13.900 ;
        RECT 105.400 13.800 106.200 13.900 ;
        RECT 102.900 12.700 103.300 12.800 ;
        RECT 99.800 12.100 100.200 12.500 ;
        RECT 101.900 12.400 103.300 12.700 ;
        RECT 103.800 12.400 104.200 12.800 ;
        RECT 101.900 12.100 102.200 12.400 ;
        RECT 104.600 12.100 105.000 12.500 ;
        RECT 99.500 11.800 100.200 12.100 ;
        RECT 99.500 11.100 100.100 11.800 ;
        RECT 101.800 11.100 102.200 12.100 ;
        RECT 104.000 11.800 105.000 12.100 ;
        RECT 104.000 11.100 104.400 11.800 ;
        RECT 106.200 11.100 106.600 13.500 ;
        RECT 107.000 12.400 107.400 13.200 ;
        RECT 107.800 11.100 108.200 14.800 ;
        RECT 110.100 14.200 110.400 15.800 ;
        RECT 111.100 15.500 113.000 15.800 ;
        RECT 111.100 14.500 111.400 15.500 ;
        RECT 109.400 13.800 110.400 14.200 ;
        RECT 110.700 14.100 111.400 14.500 ;
        RECT 111.800 14.400 112.200 15.200 ;
        RECT 112.600 14.400 113.000 15.200 ;
        RECT 110.100 13.500 110.400 13.800 ;
        RECT 110.900 13.900 111.400 14.100 ;
        RECT 110.900 13.600 113.000 13.900 ;
        RECT 110.100 13.300 110.500 13.500 ;
        RECT 110.100 13.000 110.900 13.300 ;
        RECT 110.500 11.500 110.900 13.000 ;
        RECT 112.700 12.500 113.000 13.600 ;
        RECT 112.600 11.500 113.000 12.500 ;
        RECT 113.400 12.400 113.800 13.200 ;
        RECT 114.200 11.100 114.600 15.800 ;
        RECT 115.000 17.500 115.400 19.500 ;
        RECT 115.000 15.800 115.300 17.500 ;
        RECT 117.100 16.400 117.500 19.900 ;
        RECT 117.100 16.100 117.900 16.400 ;
        RECT 115.000 15.500 116.900 15.800 ;
        RECT 115.000 14.400 115.400 15.200 ;
        RECT 115.800 14.400 116.200 15.200 ;
        RECT 116.600 14.500 116.900 15.500 ;
        RECT 116.600 14.100 117.300 14.500 ;
        RECT 117.600 14.200 117.900 16.100 ;
        RECT 118.200 14.800 118.600 15.600 ;
        RECT 119.800 15.100 120.200 15.200 ;
        RECT 120.600 15.100 121.000 19.900 ;
        RECT 121.400 17.500 121.800 19.500 ;
        RECT 121.400 15.800 121.700 17.500 ;
        RECT 123.500 16.400 123.900 19.900 ;
        RECT 123.500 16.100 124.300 16.400 ;
        RECT 121.400 15.500 123.300 15.800 ;
        RECT 119.800 14.800 121.000 15.100 ;
        RECT 116.600 13.900 117.100 14.100 ;
        RECT 115.000 13.600 117.100 13.900 ;
        RECT 117.600 13.800 118.600 14.200 ;
        RECT 115.000 12.500 115.300 13.600 ;
        RECT 117.600 13.500 117.900 13.800 ;
        RECT 117.500 13.300 117.900 13.500 ;
        RECT 117.100 13.000 117.900 13.300 ;
        RECT 115.000 11.500 115.400 12.500 ;
        RECT 117.100 12.200 117.500 13.000 ;
        RECT 119.800 12.400 120.200 13.200 ;
        RECT 116.600 11.800 117.500 12.200 ;
        RECT 117.100 11.500 117.500 11.800 ;
        RECT 120.600 11.100 121.000 14.800 ;
        RECT 121.400 14.400 121.800 15.200 ;
        RECT 122.200 14.400 122.600 15.200 ;
        RECT 123.000 14.500 123.300 15.500 ;
        RECT 123.000 14.100 123.700 14.500 ;
        RECT 124.000 14.200 124.300 16.100 ;
        RECT 126.200 15.700 126.600 19.900 ;
        RECT 128.400 18.200 128.800 19.900 ;
        RECT 127.800 17.900 128.800 18.200 ;
        RECT 130.600 17.900 131.000 19.900 ;
        RECT 132.700 17.900 133.300 19.900 ;
        RECT 127.800 17.500 128.200 17.900 ;
        RECT 130.600 17.600 130.900 17.900 ;
        RECT 129.500 17.300 131.300 17.600 ;
        RECT 132.600 17.500 133.000 17.900 ;
        RECT 129.500 17.200 129.900 17.300 ;
        RECT 130.900 17.200 131.300 17.300 ;
        RECT 127.800 16.500 128.200 16.600 ;
        RECT 130.100 16.500 130.500 16.600 ;
        RECT 127.800 16.200 130.500 16.500 ;
        RECT 130.800 16.500 131.900 16.800 ;
        RECT 130.800 15.900 131.100 16.500 ;
        RECT 131.500 16.400 131.900 16.500 ;
        RECT 132.700 16.600 133.400 17.000 ;
        RECT 132.700 16.100 133.000 16.600 ;
        RECT 128.700 15.700 131.100 15.900 ;
        RECT 126.200 15.600 131.100 15.700 ;
        RECT 131.800 15.800 133.000 16.100 ;
        RECT 124.600 14.800 125.000 15.600 ;
        RECT 126.200 15.500 129.100 15.600 ;
        RECT 126.200 15.400 129.000 15.500 ;
        RECT 129.400 15.100 129.800 15.200 ;
        RECT 127.300 14.800 129.800 15.100 ;
        RECT 127.300 14.700 127.700 14.800 ;
        RECT 128.100 14.200 128.500 14.300 ;
        RECT 131.800 14.200 132.100 15.800 ;
        RECT 135.000 15.600 135.400 19.900 ;
        RECT 133.300 15.300 135.400 15.600 ;
        RECT 133.300 15.200 133.700 15.300 ;
        RECT 134.100 14.900 134.500 15.000 ;
        RECT 132.600 14.600 134.500 14.900 ;
        RECT 132.600 14.500 133.000 14.600 ;
        RECT 123.000 13.900 123.500 14.100 ;
        RECT 121.400 13.600 123.500 13.900 ;
        RECT 124.000 13.800 125.000 14.200 ;
        RECT 126.600 13.900 132.100 14.200 ;
        RECT 126.600 13.800 127.400 13.900 ;
        RECT 121.400 12.500 121.700 13.600 ;
        RECT 124.000 13.500 124.300 13.800 ;
        RECT 123.900 13.300 124.300 13.500 ;
        RECT 123.500 13.000 124.300 13.300 ;
        RECT 121.400 11.500 121.800 12.500 ;
        RECT 123.500 12.200 123.900 13.000 ;
        RECT 123.000 11.800 123.900 12.200 ;
        RECT 123.500 11.500 123.900 11.800 ;
        RECT 126.200 11.100 126.600 13.500 ;
        RECT 128.700 12.800 129.000 13.900 ;
        RECT 131.500 13.800 131.900 13.900 ;
        RECT 135.000 13.600 135.400 15.300 ;
        RECT 133.500 13.300 135.400 13.600 ;
        RECT 133.500 13.200 133.900 13.300 ;
        RECT 135.000 13.100 135.400 13.300 ;
        RECT 136.600 15.100 137.000 19.900 ;
        RECT 139.300 16.400 139.700 19.900 ;
        RECT 141.400 17.500 141.800 19.500 ;
        RECT 138.900 16.100 139.700 16.400 ;
        RECT 138.200 15.100 138.600 15.600 ;
        RECT 136.600 14.800 138.600 15.100 ;
        RECT 135.800 13.100 136.200 13.200 ;
        RECT 135.000 12.800 136.200 13.100 ;
        RECT 127.800 12.100 128.200 12.500 ;
        RECT 128.600 12.400 129.000 12.800 ;
        RECT 129.500 12.700 129.900 12.800 ;
        RECT 129.500 12.400 130.900 12.700 ;
        RECT 130.600 12.100 130.900 12.400 ;
        RECT 132.600 12.100 133.000 12.500 ;
        RECT 127.800 11.800 128.800 12.100 ;
        RECT 128.400 11.100 128.800 11.800 ;
        RECT 130.600 11.100 131.000 12.100 ;
        RECT 132.600 11.800 133.300 12.100 ;
        RECT 132.700 11.100 133.300 11.800 ;
        RECT 135.000 11.100 135.400 12.800 ;
        RECT 135.800 12.400 136.200 12.800 ;
        RECT 136.600 11.100 137.000 14.800 ;
        RECT 138.900 14.200 139.200 16.100 ;
        RECT 141.500 15.800 141.800 17.500 ;
        RECT 145.700 19.200 146.100 19.900 ;
        RECT 145.700 18.800 146.600 19.200 ;
        RECT 145.700 16.400 146.100 18.800 ;
        RECT 147.800 17.500 148.200 19.500 ;
        RECT 139.900 15.500 141.800 15.800 ;
        RECT 145.300 16.100 146.100 16.400 ;
        RECT 139.900 14.500 140.200 15.500 ;
        RECT 138.200 13.800 139.200 14.200 ;
        RECT 139.500 14.100 140.200 14.500 ;
        RECT 140.600 14.400 141.000 15.200 ;
        RECT 141.400 15.100 141.800 15.200 ;
        RECT 143.000 15.100 143.400 15.200 ;
        RECT 141.400 14.800 143.400 15.100 ;
        RECT 144.600 14.800 145.000 15.600 ;
        RECT 141.400 14.400 141.800 14.800 ;
        RECT 145.300 14.200 145.600 16.100 ;
        RECT 147.900 15.800 148.200 17.500 ;
        RECT 146.300 15.500 148.200 15.800 ;
        RECT 148.600 17.500 149.000 19.500 ;
        RECT 148.600 15.800 148.900 17.500 ;
        RECT 150.700 16.400 151.100 19.900 ;
        RECT 150.700 16.100 151.500 16.400 ;
        RECT 148.600 15.500 150.500 15.800 ;
        RECT 146.300 14.500 146.600 15.500 ;
        RECT 138.900 13.500 139.200 13.800 ;
        RECT 139.700 13.900 140.200 14.100 ;
        RECT 139.700 13.600 141.800 13.900 ;
        RECT 144.600 13.800 145.600 14.200 ;
        RECT 145.900 14.100 146.600 14.500 ;
        RECT 147.000 14.400 147.400 15.200 ;
        RECT 147.800 14.400 148.200 15.200 ;
        RECT 148.600 14.400 149.000 15.200 ;
        RECT 149.400 14.400 149.800 15.200 ;
        RECT 150.200 14.500 150.500 15.500 ;
        RECT 138.900 13.300 139.300 13.500 ;
        RECT 138.900 13.000 139.700 13.300 ;
        RECT 139.300 11.500 139.700 13.000 ;
        RECT 141.500 12.500 141.800 13.600 ;
        RECT 145.300 13.500 145.600 13.800 ;
        RECT 146.100 13.900 146.600 14.100 ;
        RECT 150.200 14.100 150.900 14.500 ;
        RECT 151.200 14.200 151.500 16.100 ;
        RECT 153.400 15.700 153.800 19.900 ;
        RECT 155.600 18.200 156.000 19.900 ;
        RECT 155.000 17.900 156.000 18.200 ;
        RECT 157.800 17.900 158.200 19.900 ;
        RECT 159.900 17.900 160.500 19.900 ;
        RECT 155.000 17.500 155.400 17.900 ;
        RECT 157.800 17.600 158.100 17.900 ;
        RECT 156.700 17.300 158.500 17.600 ;
        RECT 159.800 17.500 160.200 17.900 ;
        RECT 156.700 17.200 157.100 17.300 ;
        RECT 158.100 17.200 158.500 17.300 ;
        RECT 155.000 16.500 155.400 16.600 ;
        RECT 157.300 16.500 157.700 16.600 ;
        RECT 155.000 16.200 157.700 16.500 ;
        RECT 158.000 16.500 159.100 16.800 ;
        RECT 158.000 15.900 158.300 16.500 ;
        RECT 158.700 16.400 159.100 16.500 ;
        RECT 159.900 16.600 160.600 17.000 ;
        RECT 159.900 16.100 160.200 16.600 ;
        RECT 155.900 15.700 158.300 15.900 ;
        RECT 153.400 15.600 158.300 15.700 ;
        RECT 159.000 15.800 160.200 16.100 ;
        RECT 151.800 15.100 152.200 15.600 ;
        RECT 153.400 15.500 156.300 15.600 ;
        RECT 153.400 15.400 156.200 15.500 ;
        RECT 152.600 15.100 153.000 15.200 ;
        RECT 156.600 15.100 157.000 15.200 ;
        RECT 151.800 14.800 153.000 15.100 ;
        RECT 154.500 14.800 157.000 15.100 ;
        RECT 158.200 15.100 158.600 15.200 ;
        RECT 159.000 15.100 159.300 15.800 ;
        RECT 162.200 15.600 162.600 19.900 ;
        RECT 160.500 15.300 162.600 15.600 ;
        RECT 163.000 17.500 163.400 19.500 ;
        RECT 165.100 19.200 165.500 19.900 ;
        RECT 164.600 18.800 165.500 19.200 ;
        RECT 163.000 15.800 163.300 17.500 ;
        RECT 165.100 16.400 165.500 18.800 ;
        RECT 165.100 16.100 165.900 16.400 ;
        RECT 163.000 15.500 164.900 15.800 ;
        RECT 160.500 15.200 160.900 15.300 ;
        RECT 158.200 14.800 159.300 15.100 ;
        RECT 161.300 14.900 161.700 15.000 ;
        RECT 154.500 14.700 154.900 14.800 ;
        RECT 155.800 14.700 156.200 14.800 ;
        RECT 155.300 14.200 155.700 14.300 ;
        RECT 159.000 14.200 159.300 14.800 ;
        RECT 159.800 14.600 161.700 14.900 ;
        RECT 159.800 14.500 160.200 14.600 ;
        RECT 150.200 13.900 150.700 14.100 ;
        RECT 146.100 13.600 148.200 13.900 ;
        RECT 145.300 13.300 145.700 13.500 ;
        RECT 145.300 13.000 146.100 13.300 ;
        RECT 141.400 11.500 141.800 12.500 ;
        RECT 145.700 11.500 146.100 13.000 ;
        RECT 147.900 12.500 148.200 13.600 ;
        RECT 147.800 11.500 148.200 12.500 ;
        RECT 148.600 13.600 150.700 13.900 ;
        RECT 151.200 13.800 152.200 14.200 ;
        RECT 153.800 13.900 159.300 14.200 ;
        RECT 153.800 13.800 154.600 13.900 ;
        RECT 148.600 12.500 148.900 13.600 ;
        RECT 151.200 13.500 151.500 13.800 ;
        RECT 151.100 13.300 151.500 13.500 ;
        RECT 150.700 13.000 151.500 13.300 ;
        RECT 148.600 11.500 149.000 12.500 ;
        RECT 150.700 11.500 151.100 13.000 ;
        RECT 153.400 11.100 153.800 13.500 ;
        RECT 155.900 12.800 156.200 13.900 ;
        RECT 158.700 13.800 159.100 13.900 ;
        RECT 162.200 13.600 162.600 15.300 ;
        RECT 163.000 14.400 163.400 15.200 ;
        RECT 163.800 14.400 164.200 15.200 ;
        RECT 164.600 14.500 164.900 15.500 ;
        RECT 164.600 14.100 165.300 14.500 ;
        RECT 165.600 14.200 165.900 16.100 ;
        RECT 166.200 14.800 166.600 15.600 ;
        RECT 164.600 13.900 165.100 14.100 ;
        RECT 160.700 13.300 162.600 13.600 ;
        RECT 160.700 13.200 161.100 13.300 ;
        RECT 155.000 12.100 155.400 12.500 ;
        RECT 155.800 12.400 156.200 12.800 ;
        RECT 156.700 12.700 157.100 12.800 ;
        RECT 156.700 12.400 158.100 12.700 ;
        RECT 157.800 12.100 158.100 12.400 ;
        RECT 159.800 12.100 160.200 12.500 ;
        RECT 155.000 11.800 156.000 12.100 ;
        RECT 155.600 11.100 156.000 11.800 ;
        RECT 157.800 11.100 158.200 12.100 ;
        RECT 159.800 11.800 160.500 12.100 ;
        RECT 159.900 11.100 160.500 11.800 ;
        RECT 162.200 11.100 162.600 13.300 ;
        RECT 163.000 13.600 165.100 13.900 ;
        RECT 165.600 13.800 166.600 14.200 ;
        RECT 163.000 12.500 163.300 13.600 ;
        RECT 165.600 13.500 165.900 13.800 ;
        RECT 165.500 13.300 165.900 13.500 ;
        RECT 167.800 13.400 168.200 14.200 ;
        RECT 165.100 13.000 165.900 13.300 ;
        RECT 168.600 13.100 169.000 19.900 ;
        RECT 169.400 15.800 169.800 16.600 ;
        RECT 170.200 16.100 170.600 19.900 ;
        RECT 171.000 16.100 171.400 16.200 ;
        RECT 170.200 15.800 171.400 16.100 ;
        RECT 171.800 16.100 172.200 16.200 ;
        RECT 172.600 16.100 173.000 19.900 ;
        RECT 171.800 15.800 173.000 16.100 ;
        RECT 163.000 11.500 163.400 12.500 ;
        RECT 165.100 11.500 165.500 13.000 ;
        RECT 168.600 12.800 169.500 13.100 ;
        RECT 169.100 11.100 169.500 12.800 ;
        RECT 170.200 11.100 170.600 15.800 ;
        RECT 171.000 12.400 171.400 13.200 ;
        RECT 171.800 12.400 172.200 13.200 ;
        RECT 172.600 11.100 173.000 15.800 ;
        RECT 173.400 11.100 173.800 19.900 ;
        RECT 176.900 16.400 177.300 19.900 ;
        RECT 179.000 17.500 179.400 19.500 ;
        RECT 176.500 16.100 177.300 16.400 ;
        RECT 175.800 14.800 176.200 15.600 ;
        RECT 176.500 14.200 176.800 16.100 ;
        RECT 179.100 15.800 179.400 17.500 ;
        RECT 177.500 15.500 179.400 15.800 ;
        RECT 177.500 14.500 177.800 15.500 ;
        RECT 175.800 13.800 176.800 14.200 ;
        RECT 177.100 14.100 177.800 14.500 ;
        RECT 178.200 14.400 178.600 15.200 ;
        RECT 179.000 14.400 179.400 15.200 ;
        RECT 176.500 13.500 176.800 13.800 ;
        RECT 177.300 13.900 177.800 14.100 ;
        RECT 177.300 13.600 179.400 13.900 ;
        RECT 176.500 13.300 176.900 13.500 ;
        RECT 174.200 12.400 174.600 13.200 ;
        RECT 176.500 13.000 177.300 13.300 ;
        RECT 176.900 12.200 177.300 13.000 ;
        RECT 179.100 12.500 179.400 13.600 ;
        RECT 176.600 11.800 177.300 12.200 ;
        RECT 176.900 11.500 177.300 11.800 ;
        RECT 179.000 11.500 179.400 12.500 ;
        RECT 0.600 7.500 1.000 9.900 ;
        RECT 2.800 9.200 3.200 9.900 ;
        RECT 2.200 8.900 3.200 9.200 ;
        RECT 5.000 8.900 5.400 9.900 ;
        RECT 7.100 9.200 7.700 9.900 ;
        RECT 7.000 8.900 7.700 9.200 ;
        RECT 2.200 8.500 2.600 8.900 ;
        RECT 5.000 8.600 5.300 8.900 ;
        RECT 3.000 8.200 3.400 8.600 ;
        RECT 3.900 8.300 5.300 8.600 ;
        RECT 7.000 8.500 7.400 8.900 ;
        RECT 3.900 8.200 4.300 8.300 ;
        RECT 1.000 7.100 1.800 7.200 ;
        RECT 3.100 7.100 3.400 8.200 ;
        RECT 7.900 7.700 8.300 7.800 ;
        RECT 9.400 7.700 9.800 9.900 ;
        RECT 7.900 7.400 9.800 7.700 ;
        RECT 10.200 7.500 10.600 9.900 ;
        RECT 12.400 9.200 12.800 9.900 ;
        RECT 11.800 8.900 12.800 9.200 ;
        RECT 14.600 8.900 15.000 9.900 ;
        RECT 16.700 9.200 17.300 9.900 ;
        RECT 16.600 8.900 17.300 9.200 ;
        RECT 11.800 8.500 12.200 8.900 ;
        RECT 14.600 8.600 14.900 8.900 ;
        RECT 12.600 8.200 13.000 8.600 ;
        RECT 13.500 8.300 14.900 8.600 ;
        RECT 16.600 8.500 17.000 8.900 ;
        RECT 13.500 8.200 13.900 8.300 ;
        RECT 4.600 7.100 5.000 7.200 ;
        RECT 5.900 7.100 6.300 7.200 ;
        RECT 1.000 6.800 6.500 7.100 ;
        RECT 2.500 6.700 2.900 6.800 ;
        RECT 1.700 6.200 2.100 6.300 ;
        RECT 3.000 6.200 3.400 6.300 ;
        RECT 1.700 5.900 4.200 6.200 ;
        RECT 3.800 5.800 4.200 5.900 ;
        RECT 0.600 5.500 3.400 5.600 ;
        RECT 0.600 5.400 3.500 5.500 ;
        RECT 0.600 5.300 5.500 5.400 ;
        RECT 0.600 1.100 1.000 5.300 ;
        RECT 3.100 5.100 5.500 5.300 ;
        RECT 2.200 4.500 4.900 4.800 ;
        RECT 2.200 4.400 2.600 4.500 ;
        RECT 4.500 4.400 4.900 4.500 ;
        RECT 5.200 4.500 5.500 5.100 ;
        RECT 6.200 5.200 6.500 6.800 ;
        RECT 7.000 6.400 7.400 6.500 ;
        RECT 7.000 6.100 8.900 6.400 ;
        RECT 8.500 6.000 8.900 6.100 ;
        RECT 7.700 5.700 8.100 5.800 ;
        RECT 9.400 5.700 9.800 7.400 ;
        RECT 10.600 7.100 11.400 7.200 ;
        RECT 12.700 7.100 13.000 8.200 ;
        RECT 17.500 7.700 17.900 7.800 ;
        RECT 19.000 7.700 19.400 9.900 ;
        RECT 17.500 7.400 19.400 7.700 ;
        RECT 14.200 7.100 14.600 7.200 ;
        RECT 15.500 7.100 15.900 7.200 ;
        RECT 10.600 6.800 16.100 7.100 ;
        RECT 12.100 6.700 12.500 6.800 ;
        RECT 11.300 6.200 11.700 6.300 ;
        RECT 12.600 6.200 13.000 6.300 ;
        RECT 11.300 5.900 13.800 6.200 ;
        RECT 13.400 5.800 13.800 5.900 ;
        RECT 7.700 5.400 9.800 5.700 ;
        RECT 6.200 4.900 7.400 5.200 ;
        RECT 5.900 4.500 6.300 4.600 ;
        RECT 5.200 4.200 6.300 4.500 ;
        RECT 7.100 4.400 7.400 4.900 ;
        RECT 7.100 4.000 7.800 4.400 ;
        RECT 3.900 3.700 4.300 3.800 ;
        RECT 5.300 3.700 5.700 3.800 ;
        RECT 2.200 3.100 2.600 3.500 ;
        RECT 3.900 3.400 5.700 3.700 ;
        RECT 5.000 3.100 5.300 3.400 ;
        RECT 7.000 3.100 7.400 3.500 ;
        RECT 2.200 2.800 3.200 3.100 ;
        RECT 2.800 1.100 3.200 2.800 ;
        RECT 5.000 1.100 5.400 3.100 ;
        RECT 7.100 1.100 7.700 3.100 ;
        RECT 9.400 1.100 9.800 5.400 ;
        RECT 10.200 5.500 13.000 5.600 ;
        RECT 10.200 5.400 13.100 5.500 ;
        RECT 10.200 5.300 15.100 5.400 ;
        RECT 10.200 1.100 10.600 5.300 ;
        RECT 12.700 5.100 15.100 5.300 ;
        RECT 11.800 4.500 14.500 4.800 ;
        RECT 11.800 4.400 12.200 4.500 ;
        RECT 14.100 4.400 14.500 4.500 ;
        RECT 14.800 4.500 15.100 5.100 ;
        RECT 15.800 5.200 16.100 6.800 ;
        RECT 16.600 6.400 17.000 6.500 ;
        RECT 16.600 6.100 18.500 6.400 ;
        RECT 18.100 6.000 18.500 6.100 ;
        RECT 17.300 5.700 17.700 5.800 ;
        RECT 19.000 5.700 19.400 7.400 ;
        RECT 21.400 7.900 21.800 9.900 ;
        RECT 23.800 8.900 24.200 9.900 ;
        RECT 22.100 8.200 22.500 8.600 ;
        RECT 20.600 6.400 21.000 7.200 ;
        RECT 19.800 6.100 20.200 6.200 ;
        RECT 21.400 6.100 21.700 7.900 ;
        RECT 22.200 7.800 22.600 8.200 ;
        RECT 23.000 7.800 23.400 8.600 ;
        RECT 22.200 7.100 22.500 7.800 ;
        RECT 23.900 7.200 24.200 8.900 ;
        RECT 25.400 7.500 25.800 9.900 ;
        RECT 27.600 9.200 28.000 9.900 ;
        RECT 27.000 8.900 28.000 9.200 ;
        RECT 29.800 8.900 30.200 9.900 ;
        RECT 31.900 9.200 32.500 9.900 ;
        RECT 31.800 8.900 32.500 9.200 ;
        RECT 27.000 8.500 27.400 8.900 ;
        RECT 29.800 8.600 30.100 8.900 ;
        RECT 27.800 8.200 28.200 8.600 ;
        RECT 28.700 8.300 30.100 8.600 ;
        RECT 31.800 8.500 32.200 8.900 ;
        RECT 28.700 8.200 29.100 8.300 ;
        RECT 23.800 7.100 24.200 7.200 ;
        RECT 22.200 6.800 24.200 7.100 ;
        RECT 25.800 7.100 26.600 7.200 ;
        RECT 27.900 7.100 28.200 8.200 ;
        RECT 32.700 7.700 33.100 7.800 ;
        RECT 34.200 7.700 34.600 9.900 ;
        RECT 32.700 7.400 34.600 7.700 ;
        RECT 36.600 7.500 37.000 9.900 ;
        RECT 38.800 9.200 39.200 9.900 ;
        RECT 38.200 8.900 39.200 9.200 ;
        RECT 41.000 8.900 41.400 9.900 ;
        RECT 43.100 9.200 43.700 9.900 ;
        RECT 43.000 8.900 43.700 9.200 ;
        RECT 38.200 8.500 38.600 8.900 ;
        RECT 41.000 8.600 41.300 8.900 ;
        RECT 39.000 8.200 39.400 8.600 ;
        RECT 39.900 8.300 41.300 8.600 ;
        RECT 43.000 8.500 43.400 8.900 ;
        RECT 39.900 8.200 40.300 8.300 ;
        RECT 29.400 7.100 29.800 7.200 ;
        RECT 30.700 7.100 31.100 7.200 ;
        RECT 25.800 6.800 31.300 7.100 ;
        RECT 22.200 6.100 22.600 6.200 ;
        RECT 19.800 5.800 20.600 6.100 ;
        RECT 21.400 5.800 22.600 6.100 ;
        RECT 17.300 5.400 19.400 5.700 ;
        RECT 20.200 5.600 20.600 5.800 ;
        RECT 15.800 4.900 17.000 5.200 ;
        RECT 15.500 4.500 15.900 4.600 ;
        RECT 14.800 4.200 15.900 4.500 ;
        RECT 16.700 4.400 17.000 4.900 ;
        RECT 16.700 4.000 17.400 4.400 ;
        RECT 13.500 3.700 13.900 3.800 ;
        RECT 14.900 3.700 15.300 3.800 ;
        RECT 11.800 3.100 12.200 3.500 ;
        RECT 13.500 3.400 15.300 3.700 ;
        RECT 14.600 3.100 14.900 3.400 ;
        RECT 16.600 3.100 17.000 3.500 ;
        RECT 11.800 2.800 12.800 3.100 ;
        RECT 12.400 1.100 12.800 2.800 ;
        RECT 14.600 1.100 15.000 3.100 ;
        RECT 16.700 1.100 17.300 3.100 ;
        RECT 19.000 1.100 19.400 5.400 ;
        RECT 22.200 5.100 22.500 5.800 ;
        RECT 23.900 5.100 24.200 6.800 ;
        RECT 27.300 6.700 27.700 6.800 ;
        RECT 26.500 6.200 26.900 6.300 ;
        RECT 27.800 6.200 28.200 6.300 ;
        RECT 24.600 5.400 25.000 6.200 ;
        RECT 26.500 5.900 29.000 6.200 ;
        RECT 28.600 5.800 29.000 5.900 ;
        RECT 25.400 5.500 28.200 5.600 ;
        RECT 25.400 5.400 28.300 5.500 ;
        RECT 25.400 5.300 30.300 5.400 ;
        RECT 19.800 4.800 21.800 5.100 ;
        RECT 19.800 1.100 20.200 4.800 ;
        RECT 21.400 1.100 21.800 4.800 ;
        RECT 22.200 1.100 22.600 5.100 ;
        RECT 23.800 4.700 24.700 5.100 ;
        RECT 24.300 1.100 24.700 4.700 ;
        RECT 25.400 1.100 25.800 5.300 ;
        RECT 27.900 5.100 30.300 5.300 ;
        RECT 27.000 4.500 29.700 4.800 ;
        RECT 27.000 4.400 27.400 4.500 ;
        RECT 29.300 4.400 29.700 4.500 ;
        RECT 30.000 4.500 30.300 5.100 ;
        RECT 31.000 5.200 31.300 6.800 ;
        RECT 31.800 6.400 32.200 6.500 ;
        RECT 31.800 6.100 33.700 6.400 ;
        RECT 33.300 6.000 33.700 6.100 ;
        RECT 32.500 5.700 32.900 5.800 ;
        RECT 34.200 5.700 34.600 7.400 ;
        RECT 37.000 7.100 37.800 7.200 ;
        RECT 39.100 7.100 39.400 8.200 ;
        RECT 45.400 8.100 45.800 9.900 ;
        RECT 47.000 8.900 47.400 9.900 ;
        RECT 46.200 8.100 46.600 8.600 ;
        RECT 47.100 8.100 47.400 8.900 ;
        RECT 48.700 8.200 49.100 8.600 ;
        RECT 48.600 8.100 49.000 8.200 ;
        RECT 45.400 7.800 46.600 8.100 ;
        RECT 47.000 7.800 49.000 8.100 ;
        RECT 49.400 7.800 49.800 9.900 ;
        RECT 43.900 7.700 44.300 7.800 ;
        RECT 45.400 7.700 45.800 7.800 ;
        RECT 43.900 7.400 45.800 7.700 ;
        RECT 41.900 7.100 42.300 7.200 ;
        RECT 37.000 6.800 42.500 7.100 ;
        RECT 38.500 6.700 38.900 6.800 ;
        RECT 37.700 6.200 38.100 6.300 ;
        RECT 37.700 6.100 40.200 6.200 ;
        RECT 41.400 6.100 41.800 6.200 ;
        RECT 37.700 5.900 41.800 6.100 ;
        RECT 39.800 5.800 41.800 5.900 ;
        RECT 32.500 5.400 34.600 5.700 ;
        RECT 31.000 4.900 32.200 5.200 ;
        RECT 30.700 4.500 31.100 4.600 ;
        RECT 30.000 4.200 31.100 4.500 ;
        RECT 31.900 4.400 32.200 4.900 ;
        RECT 31.900 4.000 32.600 4.400 ;
        RECT 28.700 3.700 29.100 3.800 ;
        RECT 30.100 3.700 30.500 3.800 ;
        RECT 27.000 3.100 27.400 3.500 ;
        RECT 28.700 3.400 30.500 3.700 ;
        RECT 29.800 3.100 30.100 3.400 ;
        RECT 31.800 3.100 32.200 3.500 ;
        RECT 27.000 2.800 28.000 3.100 ;
        RECT 27.600 1.100 28.000 2.800 ;
        RECT 29.800 1.100 30.200 3.100 ;
        RECT 31.900 1.100 32.500 3.100 ;
        RECT 34.200 1.100 34.600 5.400 ;
        RECT 36.600 5.500 39.400 5.600 ;
        RECT 36.600 5.400 39.500 5.500 ;
        RECT 36.600 5.300 41.500 5.400 ;
        RECT 36.600 1.100 37.000 5.300 ;
        RECT 39.100 5.100 41.500 5.300 ;
        RECT 38.200 4.500 40.900 4.800 ;
        RECT 38.200 4.400 38.600 4.500 ;
        RECT 40.500 4.400 40.900 4.500 ;
        RECT 41.200 4.500 41.500 5.100 ;
        RECT 42.200 5.200 42.500 6.800 ;
        RECT 43.000 6.400 43.400 6.500 ;
        RECT 43.000 6.100 44.900 6.400 ;
        RECT 44.500 6.000 44.900 6.100 ;
        RECT 43.700 5.700 44.100 5.800 ;
        RECT 45.400 5.700 45.800 7.400 ;
        RECT 47.100 7.200 47.400 7.800 ;
        RECT 47.000 6.800 47.400 7.200 ;
        RECT 43.700 5.400 45.800 5.700 ;
        RECT 42.200 4.900 43.400 5.200 ;
        RECT 41.900 4.500 42.300 4.600 ;
        RECT 41.200 4.200 42.300 4.500 ;
        RECT 43.100 4.400 43.400 4.900 ;
        RECT 43.100 4.000 43.800 4.400 ;
        RECT 39.900 3.700 40.300 3.800 ;
        RECT 41.300 3.700 41.700 3.800 ;
        RECT 38.200 3.100 38.600 3.500 ;
        RECT 39.900 3.400 41.700 3.700 ;
        RECT 41.000 3.100 41.300 3.400 ;
        RECT 43.000 3.100 43.400 3.500 ;
        RECT 38.200 2.800 39.200 3.100 ;
        RECT 38.800 1.100 39.200 2.800 ;
        RECT 41.000 1.100 41.400 3.100 ;
        RECT 43.100 1.100 43.700 3.100 ;
        RECT 45.400 1.100 45.800 5.400 ;
        RECT 47.100 5.100 47.400 6.800 ;
        RECT 47.800 5.400 48.200 6.200 ;
        RECT 48.600 6.100 49.000 6.200 ;
        RECT 49.500 6.100 49.800 7.800 ;
        RECT 51.800 7.500 52.200 9.900 ;
        RECT 54.000 9.200 54.400 9.900 ;
        RECT 53.400 8.900 54.400 9.200 ;
        RECT 56.200 8.900 56.600 9.900 ;
        RECT 58.300 9.200 58.900 9.900 ;
        RECT 58.200 8.900 58.900 9.200 ;
        RECT 53.400 8.500 53.800 8.900 ;
        RECT 56.200 8.600 56.500 8.900 ;
        RECT 54.200 8.200 54.600 8.600 ;
        RECT 55.100 8.300 56.500 8.600 ;
        RECT 58.200 8.500 58.600 8.900 ;
        RECT 55.100 8.200 55.500 8.300 ;
        RECT 50.200 6.400 50.600 7.200 ;
        RECT 52.200 7.100 53.000 7.200 ;
        RECT 54.300 7.100 54.600 8.200 ;
        RECT 59.100 7.700 59.500 7.800 ;
        RECT 60.600 7.700 61.000 9.900 ;
        RECT 59.100 7.400 61.000 7.700 ;
        RECT 57.100 7.100 57.500 7.200 ;
        RECT 52.200 6.800 57.700 7.100 ;
        RECT 53.700 6.700 54.100 6.800 ;
        RECT 52.900 6.200 53.300 6.300 ;
        RECT 51.000 6.100 51.400 6.200 ;
        RECT 48.600 5.800 49.800 6.100 ;
        RECT 50.600 5.800 51.400 6.100 ;
        RECT 52.900 5.900 55.400 6.200 ;
        RECT 55.000 5.800 55.400 5.900 ;
        RECT 48.700 5.100 49.000 5.800 ;
        RECT 50.600 5.600 51.000 5.800 ;
        RECT 51.800 5.500 54.600 5.600 ;
        RECT 51.800 5.400 54.700 5.500 ;
        RECT 51.800 5.300 56.700 5.400 ;
        RECT 47.000 4.700 47.900 5.100 ;
        RECT 47.500 1.100 47.900 4.700 ;
        RECT 48.600 1.100 49.000 5.100 ;
        RECT 49.400 4.800 51.400 5.100 ;
        RECT 49.400 1.100 49.800 4.800 ;
        RECT 51.000 1.100 51.400 4.800 ;
        RECT 51.800 1.100 52.200 5.300 ;
        RECT 54.300 5.100 56.700 5.300 ;
        RECT 53.400 4.500 56.100 4.800 ;
        RECT 53.400 4.400 53.800 4.500 ;
        RECT 55.700 4.400 56.100 4.500 ;
        RECT 56.400 4.500 56.700 5.100 ;
        RECT 57.400 5.200 57.700 6.800 ;
        RECT 58.200 6.400 58.600 6.500 ;
        RECT 58.200 6.100 60.100 6.400 ;
        RECT 59.700 6.000 60.100 6.100 ;
        RECT 58.900 5.700 59.300 5.800 ;
        RECT 60.600 5.700 61.000 7.400 ;
        RECT 58.900 5.400 61.000 5.700 ;
        RECT 57.400 4.900 58.600 5.200 ;
        RECT 57.100 4.500 57.500 4.600 ;
        RECT 56.400 4.200 57.500 4.500 ;
        RECT 58.300 4.400 58.600 4.900 ;
        RECT 58.300 4.000 59.000 4.400 ;
        RECT 55.100 3.700 55.500 3.800 ;
        RECT 56.500 3.700 56.900 3.800 ;
        RECT 53.400 3.100 53.800 3.500 ;
        RECT 55.100 3.400 56.900 3.700 ;
        RECT 56.200 3.100 56.500 3.400 ;
        RECT 58.200 3.100 58.600 3.500 ;
        RECT 53.400 2.800 54.400 3.100 ;
        RECT 54.000 1.100 54.400 2.800 ;
        RECT 56.200 1.100 56.600 3.100 ;
        RECT 58.300 1.100 58.900 3.100 ;
        RECT 60.600 1.100 61.000 5.400 ;
        RECT 62.200 7.600 62.600 9.900 ;
        RECT 63.800 7.600 64.200 9.900 ;
        RECT 62.200 7.200 64.200 7.600 ;
        RECT 65.400 7.700 65.800 9.900 ;
        RECT 67.500 9.200 68.100 9.900 ;
        RECT 67.500 8.900 68.200 9.200 ;
        RECT 69.800 8.900 70.200 9.900 ;
        RECT 72.000 9.200 72.400 9.900 ;
        RECT 72.000 8.900 73.000 9.200 ;
        RECT 67.800 8.500 68.200 8.900 ;
        RECT 69.900 8.600 70.200 8.900 ;
        RECT 69.900 8.300 71.300 8.600 ;
        RECT 70.900 8.200 71.300 8.300 ;
        RECT 71.800 8.200 72.200 8.600 ;
        RECT 72.600 8.500 73.000 8.900 ;
        RECT 66.900 7.700 67.300 7.800 ;
        RECT 65.400 7.400 67.300 7.700 ;
        RECT 62.200 5.800 62.600 7.200 ;
        RECT 62.200 5.400 64.200 5.800 ;
        RECT 62.200 1.100 62.600 5.400 ;
        RECT 63.800 1.100 64.200 5.400 ;
        RECT 65.400 5.700 65.800 7.400 ;
        RECT 68.900 7.100 69.300 7.200 ;
        RECT 71.800 7.100 72.100 8.200 ;
        RECT 74.200 7.500 74.600 9.900 ;
        RECT 75.000 7.500 75.400 9.900 ;
        RECT 77.200 9.200 77.600 9.900 ;
        RECT 76.600 8.900 77.600 9.200 ;
        RECT 79.400 8.900 79.800 9.900 ;
        RECT 81.500 9.200 82.100 9.900 ;
        RECT 81.400 8.900 82.100 9.200 ;
        RECT 76.600 8.500 77.000 8.900 ;
        RECT 79.400 8.600 79.700 8.900 ;
        RECT 77.400 8.200 77.800 8.600 ;
        RECT 78.300 8.300 79.700 8.600 ;
        RECT 81.400 8.500 81.800 8.900 ;
        RECT 78.300 8.200 78.700 8.300 ;
        RECT 73.400 7.100 74.200 7.200 ;
        RECT 75.400 7.100 76.200 7.200 ;
        RECT 77.500 7.100 77.800 8.200 ;
        RECT 83.800 8.100 84.200 9.900 ;
        RECT 84.600 8.100 85.000 8.600 ;
        RECT 83.800 7.800 85.000 8.100 ;
        RECT 82.300 7.700 82.700 7.800 ;
        RECT 83.800 7.700 84.200 7.800 ;
        RECT 82.300 7.400 84.200 7.700 ;
        RECT 78.200 7.100 78.600 7.200 ;
        RECT 80.300 7.100 80.700 7.200 ;
        RECT 68.700 6.800 80.900 7.100 ;
        RECT 67.800 6.400 68.200 6.500 ;
        RECT 66.300 6.100 68.200 6.400 ;
        RECT 66.300 6.000 66.700 6.100 ;
        RECT 67.100 5.700 67.500 5.800 ;
        RECT 65.400 5.400 67.500 5.700 ;
        RECT 65.400 1.100 65.800 5.400 ;
        RECT 68.700 5.200 69.000 6.800 ;
        RECT 72.300 6.700 72.700 6.800 ;
        RECT 76.900 6.700 77.300 6.800 ;
        RECT 71.800 6.200 72.200 6.300 ;
        RECT 73.100 6.200 73.500 6.300 ;
        RECT 71.000 5.900 73.500 6.200 ;
        RECT 76.100 6.200 76.500 6.300 ;
        RECT 76.100 5.900 78.600 6.200 ;
        RECT 71.000 5.800 71.400 5.900 ;
        RECT 78.200 5.800 78.600 5.900 ;
        RECT 71.800 5.500 74.600 5.600 ;
        RECT 71.700 5.400 74.600 5.500 ;
        RECT 67.800 4.900 69.000 5.200 ;
        RECT 69.700 5.300 74.600 5.400 ;
        RECT 69.700 5.100 72.100 5.300 ;
        RECT 67.800 4.400 68.100 4.900 ;
        RECT 67.400 4.000 68.100 4.400 ;
        RECT 68.900 4.500 69.300 4.600 ;
        RECT 69.700 4.500 70.000 5.100 ;
        RECT 68.900 4.200 70.000 4.500 ;
        RECT 70.300 4.500 73.000 4.800 ;
        RECT 70.300 4.400 70.700 4.500 ;
        RECT 72.600 4.400 73.000 4.500 ;
        RECT 69.500 3.700 69.900 3.800 ;
        RECT 70.900 3.700 71.300 3.800 ;
        RECT 67.800 3.100 68.200 3.500 ;
        RECT 69.500 3.400 71.300 3.700 ;
        RECT 69.900 3.100 70.200 3.400 ;
        RECT 72.600 3.100 73.000 3.500 ;
        RECT 67.500 1.100 68.100 3.100 ;
        RECT 69.800 1.100 70.200 3.100 ;
        RECT 72.000 2.800 73.000 3.100 ;
        RECT 72.000 1.100 72.400 2.800 ;
        RECT 74.200 1.100 74.600 5.300 ;
        RECT 75.000 5.500 77.800 5.600 ;
        RECT 75.000 5.400 77.900 5.500 ;
        RECT 75.000 5.300 79.900 5.400 ;
        RECT 75.000 1.100 75.400 5.300 ;
        RECT 77.500 5.100 79.900 5.300 ;
        RECT 76.600 4.500 79.300 4.800 ;
        RECT 76.600 4.400 77.000 4.500 ;
        RECT 78.900 4.400 79.300 4.500 ;
        RECT 79.600 4.500 79.900 5.100 ;
        RECT 80.600 5.200 80.900 6.800 ;
        RECT 81.400 6.400 81.800 6.500 ;
        RECT 81.400 6.100 83.300 6.400 ;
        RECT 82.900 6.000 83.300 6.100 ;
        RECT 82.100 5.700 82.500 5.800 ;
        RECT 83.800 5.700 84.200 7.400 ;
        RECT 82.100 5.400 84.200 5.700 ;
        RECT 80.600 4.900 81.800 5.200 ;
        RECT 80.300 4.500 80.700 4.600 ;
        RECT 79.600 4.200 80.700 4.500 ;
        RECT 81.500 4.400 81.800 4.900 ;
        RECT 81.500 4.000 82.200 4.400 ;
        RECT 78.300 3.700 78.700 3.800 ;
        RECT 79.700 3.700 80.100 3.800 ;
        RECT 76.600 3.100 77.000 3.500 ;
        RECT 78.300 3.400 80.100 3.700 ;
        RECT 79.400 3.100 79.700 3.400 ;
        RECT 81.400 3.100 81.800 3.500 ;
        RECT 76.600 2.800 77.600 3.100 ;
        RECT 77.200 1.100 77.600 2.800 ;
        RECT 79.400 1.100 79.800 3.100 ;
        RECT 81.500 1.100 82.100 3.100 ;
        RECT 83.800 1.100 84.200 5.400 ;
        RECT 85.400 6.100 85.800 9.900 ;
        RECT 88.100 8.000 88.500 9.500 ;
        RECT 90.200 8.500 90.600 9.500 ;
        RECT 87.700 7.700 88.500 8.000 ;
        RECT 87.700 7.500 88.100 7.700 ;
        RECT 87.700 7.200 88.000 7.500 ;
        RECT 90.300 7.400 90.600 8.500 ;
        RECT 86.200 7.100 86.600 7.200 ;
        RECT 87.000 7.100 88.000 7.200 ;
        RECT 86.200 6.800 88.000 7.100 ;
        RECT 88.500 7.100 90.600 7.400 ;
        RECT 93.400 7.600 93.800 9.900 ;
        RECT 95.000 7.600 95.400 9.900 ;
        RECT 93.400 7.200 95.400 7.600 ;
        RECT 96.600 7.700 97.000 9.900 ;
        RECT 98.700 9.200 99.300 9.900 ;
        RECT 98.700 8.900 99.400 9.200 ;
        RECT 101.000 8.900 101.400 9.900 ;
        RECT 103.200 9.200 103.600 9.900 ;
        RECT 103.200 8.900 104.200 9.200 ;
        RECT 99.000 8.500 99.400 8.900 ;
        RECT 101.100 8.600 101.400 8.900 ;
        RECT 101.100 8.300 102.500 8.600 ;
        RECT 102.100 8.200 102.500 8.300 ;
        RECT 103.000 8.200 103.400 8.600 ;
        RECT 103.800 8.500 104.200 8.900 ;
        RECT 98.100 7.700 98.500 7.800 ;
        RECT 96.600 7.400 98.500 7.700 ;
        RECT 88.500 6.900 89.000 7.100 ;
        RECT 87.000 6.100 87.400 6.200 ;
        RECT 85.400 5.800 87.400 6.100 ;
        RECT 85.400 1.100 85.800 5.800 ;
        RECT 87.000 5.400 87.400 5.800 ;
        RECT 87.700 4.900 88.000 6.800 ;
        RECT 88.300 6.500 89.000 6.900 ;
        RECT 88.700 5.500 89.000 6.500 ;
        RECT 89.400 5.800 89.800 6.600 ;
        RECT 90.200 5.800 90.600 6.600 ;
        RECT 92.600 6.100 93.000 6.200 ;
        RECT 93.400 6.100 93.800 7.200 ;
        RECT 92.600 5.800 93.800 6.100 ;
        RECT 88.700 5.200 90.600 5.500 ;
        RECT 87.700 4.600 88.500 4.900 ;
        RECT 88.100 1.100 88.500 4.600 ;
        RECT 90.300 3.500 90.600 5.200 ;
        RECT 90.200 1.500 90.600 3.500 ;
        RECT 93.400 5.400 95.400 5.800 ;
        RECT 93.400 1.100 93.800 5.400 ;
        RECT 95.000 1.100 95.400 5.400 ;
        RECT 96.600 5.700 97.000 7.400 ;
        RECT 100.100 7.100 100.500 7.200 ;
        RECT 103.000 7.100 103.300 8.200 ;
        RECT 105.400 7.500 105.800 9.900 ;
        RECT 106.500 9.200 106.900 9.900 ;
        RECT 106.500 8.800 107.400 9.200 ;
        RECT 106.500 8.200 106.900 8.800 ;
        RECT 106.500 7.900 107.400 8.200 ;
        RECT 104.600 7.100 105.400 7.200 ;
        RECT 99.900 6.800 105.400 7.100 ;
        RECT 99.000 6.400 99.400 6.500 ;
        RECT 97.500 6.100 99.400 6.400 ;
        RECT 97.500 6.000 97.900 6.100 ;
        RECT 98.300 5.700 98.700 5.800 ;
        RECT 96.600 5.400 98.700 5.700 ;
        RECT 96.600 1.100 97.000 5.400 ;
        RECT 99.900 5.200 100.200 6.800 ;
        RECT 103.500 6.700 103.900 6.800 ;
        RECT 103.000 6.200 103.400 6.300 ;
        RECT 104.300 6.200 104.700 6.300 ;
        RECT 102.200 5.900 104.700 6.200 ;
        RECT 102.200 5.800 102.600 5.900 ;
        RECT 103.000 5.500 105.800 5.600 ;
        RECT 102.900 5.400 105.800 5.500 ;
        RECT 99.000 4.900 100.200 5.200 ;
        RECT 100.900 5.300 105.800 5.400 ;
        RECT 100.900 5.100 103.300 5.300 ;
        RECT 99.000 4.400 99.300 4.900 ;
        RECT 98.600 4.000 99.300 4.400 ;
        RECT 100.100 4.500 100.500 4.600 ;
        RECT 100.900 4.500 101.200 5.100 ;
        RECT 100.100 4.200 101.200 4.500 ;
        RECT 101.500 4.500 104.200 4.800 ;
        RECT 101.500 4.400 101.900 4.500 ;
        RECT 103.800 4.400 104.200 4.500 ;
        RECT 100.700 3.700 101.100 3.800 ;
        RECT 102.100 3.700 102.500 3.800 ;
        RECT 99.000 3.100 99.400 3.500 ;
        RECT 100.700 3.400 102.500 3.700 ;
        RECT 101.100 3.100 101.400 3.400 ;
        RECT 103.800 3.100 104.200 3.500 ;
        RECT 98.700 1.100 99.300 3.100 ;
        RECT 101.000 1.100 101.400 3.100 ;
        RECT 103.200 2.800 104.200 3.100 ;
        RECT 103.200 1.100 103.600 2.800 ;
        RECT 105.400 1.100 105.800 5.300 ;
        RECT 107.000 1.100 107.400 7.900 ;
        RECT 108.600 7.500 109.000 9.900 ;
        RECT 110.800 9.200 111.200 9.900 ;
        RECT 110.200 8.900 111.200 9.200 ;
        RECT 113.000 8.900 113.400 9.900 ;
        RECT 115.100 9.200 115.700 9.900 ;
        RECT 115.000 8.900 115.700 9.200 ;
        RECT 110.200 8.500 110.600 8.900 ;
        RECT 113.000 8.600 113.300 8.900 ;
        RECT 111.000 8.200 111.400 8.600 ;
        RECT 111.900 8.300 113.300 8.600 ;
        RECT 115.000 8.500 115.400 8.900 ;
        RECT 111.900 8.200 112.300 8.300 ;
        RECT 109.000 7.100 109.800 7.200 ;
        RECT 111.100 7.100 111.400 8.200 ;
        RECT 115.900 7.700 116.300 7.800 ;
        RECT 117.400 7.700 117.800 9.900 ;
        RECT 115.900 7.400 117.800 7.700 ;
        RECT 111.800 7.100 112.200 7.200 ;
        RECT 113.900 7.100 114.300 7.200 ;
        RECT 109.000 6.800 114.500 7.100 ;
        RECT 110.500 6.700 110.900 6.800 ;
        RECT 109.700 6.200 110.100 6.300 ;
        RECT 109.700 6.100 112.200 6.200 ;
        RECT 112.600 6.100 113.000 6.200 ;
        RECT 109.700 5.900 113.000 6.100 ;
        RECT 111.800 5.800 113.000 5.900 ;
        RECT 108.600 5.500 111.400 5.600 ;
        RECT 108.600 5.400 111.500 5.500 ;
        RECT 108.600 5.300 113.500 5.400 ;
        RECT 108.600 1.100 109.000 5.300 ;
        RECT 111.100 5.100 113.500 5.300 ;
        RECT 110.200 4.500 112.900 4.800 ;
        RECT 110.200 4.400 110.600 4.500 ;
        RECT 112.500 4.400 112.900 4.500 ;
        RECT 113.200 4.500 113.500 5.100 ;
        RECT 114.200 5.200 114.500 6.800 ;
        RECT 115.000 6.400 115.400 6.500 ;
        RECT 115.000 6.100 116.900 6.400 ;
        RECT 116.500 6.000 116.900 6.100 ;
        RECT 115.700 5.700 116.100 5.800 ;
        RECT 117.400 5.700 117.800 7.400 ;
        RECT 115.700 5.400 117.800 5.700 ;
        RECT 114.200 4.900 115.400 5.200 ;
        RECT 113.900 4.500 114.300 4.600 ;
        RECT 113.200 4.200 114.300 4.500 ;
        RECT 115.100 4.400 115.400 4.900 ;
        RECT 115.100 4.000 115.800 4.400 ;
        RECT 111.900 3.700 112.300 3.800 ;
        RECT 113.300 3.700 113.700 3.800 ;
        RECT 110.200 3.100 110.600 3.500 ;
        RECT 111.900 3.400 113.700 3.700 ;
        RECT 113.000 3.100 113.300 3.400 ;
        RECT 115.000 3.100 115.400 3.500 ;
        RECT 110.200 2.800 111.200 3.100 ;
        RECT 110.800 1.100 111.200 2.800 ;
        RECT 113.000 1.100 113.400 3.100 ;
        RECT 115.100 1.100 115.700 3.100 ;
        RECT 117.400 1.100 117.800 5.400 ;
        RECT 119.000 7.600 119.400 9.900 ;
        RECT 120.600 7.600 121.000 9.900 ;
        RECT 123.000 8.800 123.400 9.900 ;
        RECT 119.000 7.200 121.000 7.600 ;
        RECT 123.100 7.200 123.400 8.800 ;
        RECT 119.000 5.800 119.400 7.200 ;
        RECT 123.000 6.800 123.400 7.200 ;
        RECT 121.400 6.100 121.800 6.200 ;
        RECT 120.600 5.800 121.800 6.100 ;
        RECT 119.000 5.400 121.000 5.800 ;
        RECT 119.000 1.100 119.400 5.400 ;
        RECT 120.600 1.100 121.000 5.400 ;
        RECT 123.100 5.100 123.400 6.800 ;
        RECT 123.800 6.100 124.200 6.200 ;
        RECT 124.600 6.100 125.000 9.900 ;
        RECT 126.200 7.500 126.600 9.900 ;
        RECT 128.400 9.200 128.800 9.900 ;
        RECT 127.800 8.900 128.800 9.200 ;
        RECT 130.600 8.900 131.000 9.900 ;
        RECT 132.700 9.200 133.300 9.900 ;
        RECT 132.600 8.900 133.300 9.200 ;
        RECT 127.800 8.500 128.200 8.900 ;
        RECT 130.600 8.600 130.900 8.900 ;
        RECT 128.600 8.200 129.000 8.600 ;
        RECT 129.500 8.300 130.900 8.600 ;
        RECT 132.600 8.500 133.000 8.900 ;
        RECT 129.500 8.200 129.900 8.300 ;
        RECT 126.600 7.100 127.400 7.200 ;
        RECT 128.700 7.100 129.000 8.200 ;
        RECT 133.500 7.700 133.900 7.800 ;
        RECT 135.000 7.700 135.400 9.900 ;
        RECT 137.100 9.200 137.500 9.900 ;
        RECT 136.600 8.800 137.500 9.200 ;
        RECT 137.100 8.200 137.500 8.800 ;
        RECT 133.500 7.400 135.400 7.700 ;
        RECT 136.600 7.900 137.500 8.200 ;
        RECT 131.500 7.100 131.900 7.200 ;
        RECT 135.000 7.100 135.400 7.400 ;
        RECT 135.800 7.100 136.200 7.600 ;
        RECT 126.600 6.800 132.100 7.100 ;
        RECT 128.100 6.700 128.500 6.800 ;
        RECT 123.800 5.800 125.000 6.100 ;
        RECT 127.300 6.200 127.700 6.300 ;
        RECT 127.300 5.900 129.800 6.200 ;
        RECT 129.400 5.800 129.800 5.900 ;
        RECT 123.800 5.400 124.200 5.800 ;
        RECT 123.000 4.700 123.900 5.100 ;
        RECT 123.500 1.100 123.900 4.700 ;
        RECT 124.600 1.100 125.000 5.800 ;
        RECT 126.200 5.500 129.000 5.600 ;
        RECT 126.200 5.400 129.100 5.500 ;
        RECT 126.200 5.300 131.100 5.400 ;
        RECT 126.200 1.100 126.600 5.300 ;
        RECT 128.700 5.100 131.100 5.300 ;
        RECT 127.800 4.500 130.500 4.800 ;
        RECT 127.800 4.400 128.200 4.500 ;
        RECT 130.100 4.400 130.500 4.500 ;
        RECT 130.800 4.500 131.100 5.100 ;
        RECT 131.800 5.200 132.100 6.800 ;
        RECT 135.000 6.800 136.200 7.100 ;
        RECT 132.600 6.400 133.000 6.500 ;
        RECT 132.600 6.100 134.500 6.400 ;
        RECT 134.100 6.000 134.500 6.100 ;
        RECT 133.300 5.700 133.700 5.800 ;
        RECT 135.000 5.700 135.400 6.800 ;
        RECT 133.300 5.400 135.400 5.700 ;
        RECT 131.800 4.900 133.000 5.200 ;
        RECT 131.500 4.500 131.900 4.600 ;
        RECT 130.800 4.200 131.900 4.500 ;
        RECT 132.700 4.400 133.000 4.900 ;
        RECT 132.700 4.000 133.400 4.400 ;
        RECT 129.500 3.700 129.900 3.800 ;
        RECT 130.900 3.700 131.300 3.800 ;
        RECT 127.800 3.100 128.200 3.500 ;
        RECT 129.500 3.400 131.300 3.700 ;
        RECT 130.600 3.100 130.900 3.400 ;
        RECT 132.600 3.100 133.000 3.500 ;
        RECT 127.800 2.800 128.800 3.100 ;
        RECT 128.400 1.100 128.800 2.800 ;
        RECT 130.600 1.100 131.000 3.100 ;
        RECT 132.700 1.100 133.300 3.100 ;
        RECT 135.000 1.100 135.400 5.400 ;
        RECT 136.600 1.100 137.000 7.900 ;
        RECT 138.200 7.800 138.600 8.600 ;
        RECT 139.000 6.100 139.400 9.900 ;
        RECT 143.300 8.000 143.700 9.500 ;
        RECT 145.400 8.500 145.800 9.500 ;
        RECT 142.900 7.700 143.700 8.000 ;
        RECT 142.900 7.500 143.300 7.700 ;
        RECT 142.900 7.200 143.200 7.500 ;
        RECT 145.500 7.400 145.800 8.500 ;
        RECT 139.800 7.100 140.200 7.200 ;
        RECT 142.200 7.100 143.200 7.200 ;
        RECT 139.800 6.800 143.200 7.100 ;
        RECT 143.700 7.100 145.800 7.400 ;
        RECT 146.200 8.500 146.600 9.500 ;
        RECT 146.200 7.400 146.500 8.500 ;
        RECT 148.300 8.000 148.700 9.500 ;
        RECT 148.300 7.700 149.100 8.000 ;
        RECT 148.700 7.500 149.100 7.700 ;
        RECT 151.000 7.500 151.400 9.900 ;
        RECT 153.200 9.200 153.600 9.900 ;
        RECT 152.600 8.900 153.600 9.200 ;
        RECT 155.400 8.900 155.800 9.900 ;
        RECT 157.500 9.200 158.100 9.900 ;
        RECT 157.400 8.900 158.100 9.200 ;
        RECT 152.600 8.500 153.000 8.900 ;
        RECT 155.400 8.600 155.700 8.900 ;
        RECT 153.400 8.200 153.800 8.600 ;
        RECT 154.300 8.300 155.700 8.600 ;
        RECT 157.400 8.500 157.800 8.900 ;
        RECT 154.300 8.200 154.700 8.300 ;
        RECT 146.200 7.100 148.300 7.400 ;
        RECT 143.700 6.900 144.200 7.100 ;
        RECT 142.200 6.100 142.600 6.200 ;
        RECT 139.000 5.800 142.600 6.100 ;
        RECT 137.400 4.400 137.800 5.200 ;
        RECT 139.000 1.100 139.400 5.800 ;
        RECT 142.200 5.400 142.600 5.800 ;
        RECT 142.900 4.900 143.200 6.800 ;
        RECT 143.500 6.500 144.200 6.900 ;
        RECT 147.800 6.900 148.300 7.100 ;
        RECT 148.800 7.200 149.100 7.500 ;
        RECT 148.800 7.100 149.800 7.200 ;
        RECT 150.200 7.100 150.600 7.200 ;
        RECT 143.900 5.500 144.200 6.500 ;
        RECT 144.600 5.800 145.000 6.600 ;
        RECT 145.400 6.100 145.800 6.600 ;
        RECT 146.200 6.100 146.600 6.600 ;
        RECT 145.400 5.800 146.600 6.100 ;
        RECT 147.000 5.800 147.400 6.600 ;
        RECT 147.800 6.500 148.500 6.900 ;
        RECT 148.800 6.800 150.600 7.100 ;
        RECT 151.400 7.100 152.200 7.200 ;
        RECT 153.500 7.100 153.800 8.200 ;
        RECT 158.300 7.700 158.700 7.800 ;
        RECT 159.800 7.700 160.200 9.900 ;
        RECT 158.300 7.400 160.200 7.700 ;
        RECT 160.600 7.500 161.000 9.900 ;
        RECT 162.800 9.200 163.200 9.900 ;
        RECT 162.200 8.900 163.200 9.200 ;
        RECT 165.000 8.900 165.400 9.900 ;
        RECT 167.100 9.200 167.700 9.900 ;
        RECT 167.000 8.900 167.700 9.200 ;
        RECT 162.200 8.500 162.600 8.900 ;
        RECT 165.000 8.600 165.300 8.900 ;
        RECT 163.000 8.200 163.400 8.600 ;
        RECT 163.900 8.300 165.300 8.600 ;
        RECT 167.000 8.500 167.400 8.900 ;
        RECT 163.900 8.200 164.300 8.300 ;
        RECT 154.200 7.100 154.600 7.200 ;
        RECT 156.300 7.100 156.700 7.200 ;
        RECT 151.400 6.800 156.900 7.100 ;
        RECT 147.800 5.500 148.100 6.500 ;
        RECT 143.900 5.200 145.800 5.500 ;
        RECT 142.900 4.600 143.700 4.900 ;
        RECT 143.300 1.100 143.700 4.600 ;
        RECT 145.500 3.500 145.800 5.200 ;
        RECT 145.400 1.500 145.800 3.500 ;
        RECT 146.200 5.200 148.100 5.500 ;
        RECT 146.200 3.500 146.500 5.200 ;
        RECT 148.800 4.900 149.100 6.800 ;
        RECT 152.900 6.700 153.300 6.800 ;
        RECT 152.100 6.200 152.500 6.300 ;
        RECT 153.400 6.200 153.800 6.300 ;
        RECT 149.400 5.400 149.800 6.200 ;
        RECT 152.100 5.900 154.600 6.200 ;
        RECT 154.200 5.800 154.600 5.900 ;
        RECT 151.000 5.500 153.800 5.600 ;
        RECT 151.000 5.400 153.900 5.500 ;
        RECT 148.300 4.600 149.100 4.900 ;
        RECT 151.000 5.300 155.900 5.400 ;
        RECT 146.200 1.500 146.600 3.500 ;
        RECT 148.300 1.100 148.700 4.600 ;
        RECT 151.000 1.100 151.400 5.300 ;
        RECT 153.500 5.100 155.900 5.300 ;
        RECT 152.600 4.500 155.300 4.800 ;
        RECT 152.600 4.400 153.000 4.500 ;
        RECT 154.900 4.400 155.300 4.500 ;
        RECT 155.600 4.500 155.900 5.100 ;
        RECT 156.600 5.200 156.900 6.800 ;
        RECT 157.400 6.400 157.800 6.500 ;
        RECT 157.400 6.100 159.300 6.400 ;
        RECT 158.900 6.000 159.300 6.100 ;
        RECT 158.100 5.700 158.500 5.800 ;
        RECT 159.800 5.700 160.200 7.400 ;
        RECT 161.000 7.100 161.800 7.200 ;
        RECT 163.100 7.100 163.400 8.200 ;
        RECT 167.900 7.700 168.300 7.800 ;
        RECT 169.400 7.700 169.800 9.900 ;
        RECT 167.900 7.400 169.800 7.700 ;
        RECT 170.200 7.500 170.600 9.900 ;
        RECT 172.400 9.200 172.800 9.900 ;
        RECT 171.800 8.900 172.800 9.200 ;
        RECT 174.600 8.900 175.000 9.900 ;
        RECT 176.700 9.200 177.300 9.900 ;
        RECT 176.600 8.900 177.300 9.200 ;
        RECT 171.800 8.500 172.200 8.900 ;
        RECT 174.600 8.600 174.900 8.900 ;
        RECT 172.600 8.200 173.000 8.600 ;
        RECT 173.500 8.300 174.900 8.600 ;
        RECT 176.600 8.500 177.000 8.900 ;
        RECT 173.500 8.200 173.900 8.300 ;
        RECT 165.900 7.100 166.300 7.200 ;
        RECT 161.000 6.800 166.500 7.100 ;
        RECT 162.500 6.700 162.900 6.800 ;
        RECT 161.700 6.200 162.100 6.300 ;
        RECT 161.700 5.900 164.200 6.200 ;
        RECT 163.800 5.800 164.200 5.900 ;
        RECT 158.100 5.400 160.200 5.700 ;
        RECT 156.600 4.900 157.800 5.200 ;
        RECT 156.300 4.500 156.700 4.600 ;
        RECT 155.600 4.200 156.700 4.500 ;
        RECT 157.500 4.400 157.800 4.900 ;
        RECT 157.500 4.000 158.200 4.400 ;
        RECT 154.300 3.700 154.700 3.800 ;
        RECT 155.700 3.700 156.100 3.800 ;
        RECT 152.600 3.100 153.000 3.500 ;
        RECT 154.300 3.400 156.100 3.700 ;
        RECT 155.400 3.100 155.700 3.400 ;
        RECT 157.400 3.100 157.800 3.500 ;
        RECT 152.600 2.800 153.600 3.100 ;
        RECT 153.200 1.100 153.600 2.800 ;
        RECT 155.400 1.100 155.800 3.100 ;
        RECT 157.500 1.100 158.100 3.100 ;
        RECT 159.800 1.100 160.200 5.400 ;
        RECT 160.600 5.500 163.400 5.600 ;
        RECT 160.600 5.400 163.500 5.500 ;
        RECT 160.600 5.300 165.500 5.400 ;
        RECT 160.600 1.100 161.000 5.300 ;
        RECT 163.100 5.100 165.500 5.300 ;
        RECT 162.200 4.500 164.900 4.800 ;
        RECT 162.200 4.400 162.600 4.500 ;
        RECT 164.500 4.400 164.900 4.500 ;
        RECT 165.200 4.500 165.500 5.100 ;
        RECT 166.200 5.200 166.500 6.800 ;
        RECT 167.000 6.400 167.400 6.500 ;
        RECT 167.000 6.100 168.900 6.400 ;
        RECT 168.500 6.000 168.900 6.100 ;
        RECT 167.700 5.700 168.100 5.800 ;
        RECT 169.400 5.700 169.800 7.400 ;
        RECT 170.600 7.100 171.400 7.200 ;
        RECT 172.700 7.100 173.000 8.200 ;
        RECT 177.500 7.700 177.900 7.800 ;
        RECT 179.000 7.700 179.400 9.900 ;
        RECT 177.500 7.400 179.400 7.700 ;
        RECT 175.500 7.100 175.900 7.200 ;
        RECT 170.600 6.800 176.100 7.100 ;
        RECT 172.100 6.700 172.500 6.800 ;
        RECT 171.300 6.200 171.700 6.300 ;
        RECT 172.600 6.200 173.000 6.300 ;
        RECT 171.300 5.900 173.800 6.200 ;
        RECT 173.400 5.800 173.800 5.900 ;
        RECT 167.700 5.400 169.800 5.700 ;
        RECT 166.200 4.900 167.400 5.200 ;
        RECT 165.900 4.500 166.300 4.600 ;
        RECT 165.200 4.200 166.300 4.500 ;
        RECT 167.100 4.400 167.400 4.900 ;
        RECT 167.100 4.000 167.800 4.400 ;
        RECT 163.900 3.700 164.300 3.800 ;
        RECT 165.300 3.700 165.700 3.800 ;
        RECT 162.200 3.100 162.600 3.500 ;
        RECT 163.900 3.400 165.700 3.700 ;
        RECT 165.000 3.100 165.300 3.400 ;
        RECT 167.000 3.100 167.400 3.500 ;
        RECT 162.200 2.800 163.200 3.100 ;
        RECT 162.800 1.100 163.200 2.800 ;
        RECT 165.000 1.100 165.400 3.100 ;
        RECT 167.100 1.100 167.700 3.100 ;
        RECT 169.400 1.100 169.800 5.400 ;
        RECT 170.200 5.500 173.000 5.600 ;
        RECT 170.200 5.400 173.100 5.500 ;
        RECT 170.200 5.300 175.100 5.400 ;
        RECT 170.200 1.100 170.600 5.300 ;
        RECT 172.700 5.100 175.100 5.300 ;
        RECT 171.800 4.500 174.500 4.800 ;
        RECT 171.800 4.400 172.200 4.500 ;
        RECT 174.100 4.400 174.500 4.500 ;
        RECT 174.800 4.500 175.100 5.100 ;
        RECT 175.800 5.200 176.100 6.800 ;
        RECT 176.600 6.400 177.000 6.500 ;
        RECT 176.600 6.100 178.500 6.400 ;
        RECT 178.100 6.000 178.500 6.100 ;
        RECT 177.300 5.700 177.700 5.800 ;
        RECT 179.000 5.700 179.400 7.400 ;
        RECT 177.300 5.400 179.400 5.700 ;
        RECT 175.800 4.900 177.000 5.200 ;
        RECT 175.500 4.500 175.900 4.600 ;
        RECT 174.800 4.200 175.900 4.500 ;
        RECT 176.700 4.400 177.000 4.900 ;
        RECT 176.700 4.000 177.400 4.400 ;
        RECT 173.500 3.700 173.900 3.800 ;
        RECT 174.900 3.700 175.300 3.800 ;
        RECT 171.800 3.100 172.200 3.500 ;
        RECT 173.500 3.400 175.300 3.700 ;
        RECT 174.600 3.100 174.900 3.400 ;
        RECT 176.600 3.100 177.000 3.500 ;
        RECT 171.800 2.800 172.800 3.100 ;
        RECT 172.400 1.100 172.800 2.800 ;
        RECT 174.600 1.100 175.000 3.100 ;
        RECT 176.700 1.100 177.300 3.100 ;
        RECT 179.000 1.100 179.400 5.400 ;
      LAYER via1 ;
        RECT 15.800 168.800 16.200 169.200 ;
        RECT 9.400 165.900 9.800 166.300 ;
        RECT 3.800 164.800 4.200 165.200 ;
        RECT 7.000 165.100 7.400 165.500 ;
        RECT 20.600 165.800 21.000 166.200 ;
        RECT 16.600 165.100 17.000 165.500 ;
        RECT 25.400 161.800 25.800 162.200 ;
        RECT 34.200 166.800 34.600 167.200 ;
        RECT 28.600 166.100 29.000 166.500 ;
        RECT 32.600 165.900 33.000 166.300 ;
        RECT 41.400 166.800 41.800 167.200 ;
        RECT 35.000 165.100 35.400 165.500 ;
        RECT 26.200 161.800 26.600 162.200 ;
        RECT 52.600 168.800 53.000 169.200 ;
        RECT 46.200 165.900 46.600 166.300 ;
        RECT 43.800 165.100 44.200 165.500 ;
        RECT 61.400 166.800 61.800 167.200 ;
        RECT 60.600 165.100 61.000 165.500 ;
        RECT 91.800 166.800 92.200 167.200 ;
        RECT 88.600 165.800 89.000 166.200 ;
        RECT 67.800 163.800 68.200 164.200 ;
        RECT 69.400 161.800 69.800 162.200 ;
        RECT 72.600 161.800 73.000 162.200 ;
        RECT 83.800 161.800 84.200 162.200 ;
        RECT 91.000 165.100 91.400 165.500 ;
        RECT 104.600 166.800 105.000 167.200 ;
        RECT 99.800 161.800 100.200 162.200 ;
        RECT 112.600 166.800 113.000 167.200 ;
        RECT 109.400 166.100 109.800 166.500 ;
        RECT 115.800 165.100 116.200 165.500 ;
        RECT 107.000 161.800 107.400 162.200 ;
        RECT 125.400 167.800 125.800 168.200 ;
        RECT 126.200 167.100 126.600 167.500 ;
        RECT 117.400 161.800 117.800 162.200 ;
        RECT 123.000 163.400 123.400 163.800 ;
        RECT 124.600 163.100 125.000 163.500 ;
        RECT 122.200 162.100 122.600 162.500 ;
        RECT 123.000 162.100 123.400 162.500 ;
        RECT 123.800 162.100 124.200 162.500 ;
        RECT 126.200 163.100 126.600 163.500 ;
        RECT 127.800 163.100 128.200 163.500 ;
        RECT 139.800 166.500 140.200 166.900 ;
        RECT 144.600 166.300 145.000 166.700 ;
        RECT 156.600 166.800 157.000 167.200 ;
        RECT 140.600 164.400 141.000 164.800 ;
        RECT 143.000 163.800 143.400 164.200 ;
        RECT 128.600 162.100 129.000 162.500 ;
        RECT 129.400 162.100 129.800 162.500 ;
        RECT 141.400 163.100 141.800 163.500 ;
        RECT 139.800 162.100 140.200 162.500 ;
        RECT 140.600 162.100 141.000 162.500 ;
        RECT 143.000 163.100 143.400 163.500 ;
        RECT 144.600 163.100 145.000 163.500 ;
        RECT 145.400 162.100 145.800 162.500 ;
        RECT 146.200 162.100 146.600 162.500 ;
        RECT 147.000 162.100 147.400 162.500 ;
        RECT 151.800 161.800 152.200 162.200 ;
        RECT 155.800 165.100 156.200 165.500 ;
        RECT 164.600 161.800 165.000 162.200 ;
        RECT 168.600 165.800 169.000 166.200 ;
        RECT 173.400 165.800 173.800 166.200 ;
        RECT 167.800 161.800 168.200 162.200 ;
        RECT 172.600 161.800 173.000 162.200 ;
        RECT 10.200 156.800 10.600 157.200 ;
        RECT 3.800 154.800 4.200 155.200 ;
        RECT 0.600 153.100 1.000 153.500 ;
        RECT 10.200 152.800 10.600 153.200 ;
        RECT 15.000 154.800 15.400 155.200 ;
        RECT 15.800 154.800 16.200 155.200 ;
        RECT 16.600 153.800 17.000 154.200 ;
        RECT 19.000 154.800 19.400 155.200 ;
        RECT 19.800 154.800 20.200 155.200 ;
        RECT 18.200 151.800 18.600 152.200 ;
        RECT 25.400 153.800 25.800 154.200 ;
        RECT 28.600 158.800 29.000 159.200 ;
        RECT 39.800 154.800 40.200 155.200 ;
        RECT 27.000 151.800 27.400 152.200 ;
        RECT 36.600 153.100 37.000 153.500 ;
        RECT 51.800 154.800 52.200 155.200 ;
        RECT 52.600 154.800 53.000 155.200 ;
        RECT 45.400 151.800 45.800 152.200 ;
        RECT 49.400 151.800 49.800 152.200 ;
        RECT 60.600 154.800 61.000 155.200 ;
        RECT 61.400 154.800 61.800 155.200 ;
        RECT 64.600 153.800 65.000 154.200 ;
        RECT 74.200 156.200 74.600 156.600 ;
        RECT 75.800 155.500 76.200 155.900 ;
        RECT 75.800 153.100 76.200 153.500 ;
        RECT 80.600 153.800 81.000 154.200 ;
        RECT 79.800 153.100 80.200 153.500 ;
        RECT 91.000 154.800 91.400 155.200 ;
        RECT 91.800 154.800 92.200 155.200 ;
        RECT 88.600 151.800 89.000 152.200 ;
        RECT 101.400 156.800 101.800 157.200 ;
        RECT 96.600 152.800 97.000 153.200 ;
        RECT 97.400 152.800 97.800 153.200 ;
        RECT 102.200 154.800 102.600 155.200 ;
        RECT 103.000 154.800 103.400 155.200 ;
        RECT 111.000 156.200 111.400 156.600 ;
        RECT 112.600 155.500 113.000 155.900 ;
        RECT 120.600 156.200 121.000 156.600 ;
        RECT 122.200 155.500 122.600 155.900 ;
        RECT 110.200 152.800 110.600 153.200 ;
        RECT 103.800 151.800 104.200 152.200 ;
        RECT 112.600 153.100 113.000 153.500 ;
        RECT 122.200 153.100 122.600 153.500 ;
        RECT 113.400 151.800 113.800 152.200 ;
        RECT 123.000 152.800 123.400 153.200 ;
        RECT 127.800 154.800 128.200 155.200 ;
        RECT 128.600 154.800 129.000 155.200 ;
        RECT 129.400 154.800 129.800 155.200 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 133.400 153.800 133.800 154.200 ;
        RECT 135.000 152.800 135.400 153.200 ;
        RECT 137.400 153.100 137.800 153.500 ;
        RECT 139.800 152.800 140.200 153.200 ;
        RECT 146.200 151.800 146.600 152.200 ;
        RECT 154.200 152.800 154.600 153.200 ;
        RECT 152.600 151.800 153.000 152.200 ;
        RECT 155.000 151.800 155.400 152.200 ;
        RECT 164.600 157.500 165.000 157.900 ;
        RECT 163.000 156.800 163.400 157.200 ;
        RECT 165.400 156.200 165.800 156.600 ;
        RECT 159.800 154.100 160.200 154.500 ;
        RECT 164.600 154.300 165.000 154.700 ;
        RECT 162.200 153.800 162.600 154.200 ;
        RECT 159.800 152.100 160.200 152.500 ;
        RECT 160.600 152.100 161.000 152.500 ;
        RECT 161.400 152.100 161.800 152.500 ;
        RECT 163.000 152.100 163.400 152.500 ;
        RECT 164.600 152.100 165.000 152.500 ;
        RECT 165.400 152.100 165.800 152.500 ;
        RECT 166.200 152.100 166.600 152.500 ;
        RECT 167.000 152.100 167.400 152.500 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 171.800 151.800 172.200 152.200 ;
        RECT 177.400 154.800 177.800 155.200 ;
        RECT 176.600 152.800 177.000 153.200 ;
        RECT 175.800 151.800 176.200 152.200 ;
        RECT 9.400 148.800 9.800 149.200 ;
        RECT 0.600 145.100 1.000 145.500 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 14.200 146.800 14.600 147.200 ;
        RECT 15.000 145.800 15.400 146.200 ;
        RECT 20.600 147.800 21.000 148.200 ;
        RECT 17.400 144.800 17.800 145.200 ;
        RECT 25.400 146.800 25.800 147.200 ;
        RECT 35.800 146.800 36.200 147.200 ;
        RECT 39.800 146.800 40.200 147.200 ;
        RECT 30.200 146.100 30.600 146.500 ;
        RECT 42.200 145.800 42.600 146.200 ;
        RECT 36.600 145.100 37.000 145.500 ;
        RECT 27.800 141.800 28.200 142.200 ;
        RECT 41.400 144.800 41.800 145.200 ;
        RECT 55.800 148.800 56.200 149.200 ;
        RECT 49.400 145.900 49.800 146.300 ;
        RECT 46.200 144.800 46.600 145.200 ;
        RECT 47.000 145.100 47.400 145.500 ;
        RECT 45.400 141.800 45.800 142.200 ;
        RECT 67.000 146.800 67.400 147.200 ;
        RECT 71.000 146.100 71.400 146.500 ;
        RECT 59.000 143.800 59.400 144.200 ;
        RECT 58.200 141.800 58.600 142.200 ;
        RECT 61.400 144.800 61.800 145.200 ;
        RECT 75.000 145.900 75.400 146.300 ;
        RECT 78.200 145.800 78.600 146.200 ;
        RECT 77.400 145.100 77.800 145.500 ;
        RECT 84.600 146.800 85.000 147.200 ;
        RECT 93.400 146.800 93.800 147.200 ;
        RECT 99.000 147.800 99.400 148.200 ;
        RECT 91.000 146.100 91.400 146.500 ;
        RECT 97.400 145.100 97.800 145.500 ;
        RECT 88.600 141.800 89.000 142.200 ;
        RECT 98.200 144.800 98.600 145.200 ;
        RECT 104.600 146.800 105.000 147.200 ;
        RECT 105.400 146.800 105.800 147.200 ;
        RECT 100.600 145.800 101.000 146.200 ;
        RECT 104.600 145.800 105.000 146.200 ;
        RECT 108.600 145.800 109.000 146.200 ;
        RECT 107.000 141.800 107.400 142.200 ;
        RECT 117.400 144.800 117.800 145.200 ;
        RECT 131.000 146.800 131.400 147.200 ;
        RECT 123.800 146.100 124.200 146.500 ;
        RECT 131.800 145.800 132.200 146.200 ;
        RECT 130.200 145.100 130.600 145.500 ;
        RECT 121.400 141.800 121.800 142.200 ;
        RECT 136.600 145.800 137.000 146.200 ;
        RECT 132.600 144.800 133.000 145.200 ;
        RECT 150.200 148.800 150.600 149.200 ;
        RECT 147.000 146.800 147.400 147.200 ;
        RECT 149.400 146.800 149.800 147.200 ;
        RECT 141.400 146.100 141.800 146.500 ;
        RECT 147.800 145.100 148.200 145.500 ;
        RECT 158.200 148.800 158.600 149.200 ;
        RECT 157.400 146.800 157.800 147.200 ;
        RECT 154.200 145.800 154.600 146.200 ;
        RECT 159.800 145.800 160.200 146.200 ;
        RECT 166.200 146.500 166.600 146.900 ;
        RECT 171.000 146.300 171.400 146.700 ;
        RECT 167.000 144.400 167.400 144.800 ;
        RECT 169.400 143.800 169.800 144.200 ;
        RECT 167.800 143.100 168.200 143.500 ;
        RECT 166.200 142.100 166.600 142.500 ;
        RECT 167.000 142.100 167.400 142.500 ;
        RECT 169.400 143.100 169.800 143.500 ;
        RECT 171.000 143.100 171.400 143.500 ;
        RECT 171.800 142.100 172.200 142.500 ;
        RECT 172.600 142.100 173.000 142.500 ;
        RECT 173.400 142.100 173.800 142.500 ;
        RECT 178.200 141.800 178.600 142.200 ;
        RECT 19.000 136.800 19.400 137.200 ;
        RECT 0.600 133.100 1.000 133.500 ;
        RECT 13.400 134.800 13.800 135.200 ;
        RECT 11.000 133.800 11.400 134.200 ;
        RECT 9.400 131.800 9.800 132.200 ;
        RECT 10.200 133.100 10.600 133.500 ;
        RECT 15.800 133.800 16.200 134.200 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 20.600 134.800 21.000 135.200 ;
        RECT 28.600 138.800 29.000 139.200 ;
        RECT 25.400 132.800 25.800 133.200 ;
        RECT 29.400 133.800 29.800 134.200 ;
        RECT 33.400 136.800 33.800 137.200 ;
        RECT 36.600 136.800 37.000 137.200 ;
        RECT 31.800 135.800 32.200 136.200 ;
        RECT 43.800 134.800 44.200 135.200 ;
        RECT 57.400 138.800 57.800 139.200 ;
        RECT 56.600 136.800 57.000 137.200 ;
        RECT 38.200 132.800 38.600 133.200 ;
        RECT 39.800 133.100 40.200 133.500 ;
        RECT 48.600 131.800 49.000 132.200 ;
        RECT 55.000 135.800 55.400 136.200 ;
        RECT 51.000 132.800 51.400 133.200 ;
        RECT 58.200 133.800 58.600 134.200 ;
        RECT 62.200 136.800 62.600 137.200 ;
        RECT 60.600 135.800 61.000 136.200 ;
        RECT 63.800 133.800 64.200 134.200 ;
        RECT 67.800 133.800 68.200 134.200 ;
        RECT 68.600 133.800 69.000 134.200 ;
        RECT 59.800 131.800 60.200 132.200 ;
        RECT 75.000 138.800 75.400 139.200 ;
        RECT 67.000 131.800 67.400 132.200 ;
        RECT 70.200 131.800 70.600 132.200 ;
        RECT 72.600 134.800 73.000 135.200 ;
        RECT 73.400 134.800 73.800 135.200 ;
        RECT 71.800 132.800 72.200 133.200 ;
        RECT 79.000 133.800 79.400 134.200 ;
        RECT 81.400 133.800 81.800 134.200 ;
        RECT 103.800 136.200 104.200 136.600 ;
        RECT 105.400 135.500 105.800 135.900 ;
        RECT 110.200 134.800 110.600 135.200 ;
        RECT 80.600 131.800 81.000 132.200 ;
        RECT 88.600 131.800 89.000 132.200 ;
        RECT 94.200 131.800 94.600 132.200 ;
        RECT 105.400 133.100 105.800 133.500 ;
        RECT 96.600 131.800 97.000 132.200 ;
        RECT 110.200 132.800 110.600 133.200 ;
        RECT 115.000 134.800 115.400 135.200 ;
        RECT 115.800 134.800 116.200 135.200 ;
        RECT 119.800 134.800 120.200 135.200 ;
        RECT 116.600 133.100 117.000 133.500 ;
        RECT 131.000 134.800 131.400 135.200 ;
        RECT 131.800 134.800 132.200 135.200 ;
        RECT 134.200 134.800 134.600 135.200 ;
        RECT 135.800 134.800 136.200 135.200 ;
        RECT 137.400 134.800 137.800 135.200 ;
        RECT 146.200 136.200 146.600 136.600 ;
        RECT 147.800 135.500 148.200 135.900 ;
        RECT 147.800 133.100 148.200 133.500 ;
        RECT 151.000 133.800 151.400 134.200 ;
        RECT 139.000 131.800 139.400 132.200 ;
        RECT 148.600 131.800 149.000 132.200 ;
        RECT 151.800 132.800 152.200 133.200 ;
        RECT 163.000 138.800 163.400 139.200 ;
        RECT 156.600 134.800 157.000 135.200 ;
        RECT 157.400 134.800 157.800 135.200 ;
        RECT 159.800 132.800 160.200 133.200 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 167.800 134.800 168.200 135.200 ;
        RECT 168.600 134.800 169.000 135.200 ;
        RECT 167.000 133.800 167.400 134.200 ;
        RECT 172.600 134.800 173.000 135.200 ;
        RECT 173.400 134.800 173.800 135.200 ;
        RECT 179.800 132.800 180.200 133.200 ;
        RECT 3.000 128.800 3.400 129.200 ;
        RECT 1.400 125.800 1.800 126.200 ;
        RECT 6.200 125.800 6.600 126.200 ;
        RECT 11.000 126.800 11.400 127.200 ;
        RECT 22.200 128.800 22.600 129.200 ;
        RECT 15.800 125.900 16.200 126.300 ;
        RECT 13.400 125.100 13.800 125.500 ;
        RECT 35.000 128.800 35.400 129.200 ;
        RECT 27.000 126.800 27.400 127.200 ;
        RECT 26.200 125.100 26.600 125.500 ;
        RECT 25.400 121.800 25.800 122.200 ;
        RECT 59.000 128.800 59.400 129.200 ;
        RECT 51.000 126.800 51.400 127.200 ;
        RECT 50.200 125.100 50.600 125.500 ;
        RECT 60.600 127.800 61.000 128.200 ;
        RECT 79.800 128.800 80.200 129.200 ;
        RECT 61.400 125.800 61.800 126.200 ;
        RECT 67.800 125.800 68.200 126.200 ;
        RECT 85.400 126.800 85.800 127.200 ;
        RECT 86.200 125.800 86.600 126.200 ;
        RECT 82.200 125.100 82.600 125.500 ;
        RECT 71.800 121.800 72.200 122.200 ;
        RECT 75.000 121.800 75.400 122.200 ;
        RECT 103.800 128.800 104.200 129.200 ;
        RECT 93.400 123.800 93.800 124.200 ;
        RECT 107.800 128.800 108.200 129.200 ;
        RECT 103.000 126.800 103.400 127.200 ;
        RECT 99.800 124.800 100.200 125.200 ;
        RECT 105.400 125.800 105.800 126.200 ;
        RECT 117.400 128.800 117.800 129.200 ;
        RECT 115.800 126.800 116.200 127.200 ;
        RECT 110.200 126.100 110.600 126.500 ;
        RECT 119.800 126.100 120.200 126.500 ;
        RECT 116.600 125.100 117.000 125.500 ;
        RECT 123.800 125.900 124.200 126.300 ;
        RECT 126.200 125.100 126.600 125.500 ;
        RECT 133.400 126.800 133.800 127.200 ;
        RECT 142.200 128.800 142.600 129.200 ;
        RECT 139.000 127.800 139.400 128.200 ;
        RECT 147.800 128.800 148.200 129.200 ;
        RECT 150.200 128.800 150.600 129.200 ;
        RECT 131.800 125.800 132.200 126.200 ;
        RECT 149.400 127.800 149.800 128.200 ;
        RECT 148.600 126.800 149.000 127.200 ;
        RECT 147.000 125.800 147.400 126.200 ;
        RECT 155.800 126.800 156.200 127.200 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 152.600 126.100 153.000 126.500 ;
        RECT 159.000 125.100 159.400 125.500 ;
        RECT 175.000 126.800 175.400 127.200 ;
        RECT 167.000 125.800 167.400 126.200 ;
        RECT 168.600 125.800 169.000 126.200 ;
        RECT 166.200 124.800 166.600 125.200 ;
        RECT 173.400 125.900 173.800 126.300 ;
        RECT 171.000 125.100 171.400 125.500 ;
        RECT 179.800 121.800 180.200 122.200 ;
        RECT 3.000 116.800 3.400 117.200 ;
        RECT 3.800 114.800 4.200 115.200 ;
        RECT 4.600 114.800 5.000 115.200 ;
        RECT 15.800 116.800 16.200 117.200 ;
        RECT 6.200 114.800 6.600 115.200 ;
        RECT 6.200 112.800 6.600 113.200 ;
        RECT 7.000 113.100 7.400 113.500 ;
        RECT 25.400 114.800 25.800 115.200 ;
        RECT 39.800 118.800 40.200 119.200 ;
        RECT 18.200 111.800 18.600 112.200 ;
        RECT 21.400 112.800 21.800 113.200 ;
        RECT 22.200 113.100 22.600 113.500 ;
        RECT 24.600 112.800 25.000 113.200 ;
        RECT 31.000 111.800 31.400 112.200 ;
        RECT 33.400 112.800 33.800 113.200 ;
        RECT 36.600 112.800 37.000 113.200 ;
        RECT 43.800 116.800 44.200 117.200 ;
        RECT 41.400 114.800 41.800 115.200 ;
        RECT 42.200 114.800 42.600 115.200 ;
        RECT 56.600 116.800 57.000 117.200 ;
        RECT 55.000 115.800 55.400 116.200 ;
        RECT 47.000 112.800 47.400 113.200 ;
        RECT 47.800 113.100 48.200 113.500 ;
        RECT 64.600 116.200 65.000 116.600 ;
        RECT 66.200 115.500 66.600 115.900 ;
        RECT 66.200 113.100 66.600 113.500 ;
        RECT 57.400 111.800 57.800 112.200 ;
        RECT 67.000 112.800 67.400 113.200 ;
        RECT 81.400 118.800 81.800 119.200 ;
        RECT 80.600 116.800 81.000 117.200 ;
        RECT 71.800 114.800 72.200 115.200 ;
        RECT 72.600 114.800 73.000 115.200 ;
        RECT 81.400 114.800 81.800 115.200 ;
        RECT 71.000 111.800 71.400 112.200 ;
        RECT 79.000 111.800 79.400 112.200 ;
        RECT 85.400 114.800 85.800 115.200 ;
        RECT 86.200 114.800 86.600 115.200 ;
        RECT 84.600 113.800 85.000 114.200 ;
        RECT 95.800 117.800 96.200 118.200 ;
        RECT 91.000 113.800 91.400 114.200 ;
        RECT 92.600 112.800 93.000 113.200 ;
        RECT 99.800 116.800 100.200 117.200 ;
        RECT 99.000 113.800 99.400 114.200 ;
        RECT 107.000 116.200 107.400 116.600 ;
        RECT 108.600 115.500 109.000 115.900 ;
        RECT 112.600 115.800 113.000 116.200 ;
        RECT 108.600 113.100 109.000 113.500 ;
        RECT 109.400 112.800 109.800 113.200 ;
        RECT 114.200 114.800 114.600 115.200 ;
        RECT 115.000 114.800 115.400 115.200 ;
        RECT 123.000 116.200 123.400 116.600 ;
        RECT 124.600 115.500 125.000 115.900 ;
        RECT 139.000 116.800 139.400 117.200 ;
        RECT 132.600 114.800 133.000 115.200 ;
        RECT 133.400 114.800 133.800 115.200 ;
        RECT 124.600 113.100 125.000 113.500 ;
        RECT 115.800 111.800 116.200 112.200 ;
        RECT 126.200 111.800 126.600 112.200 ;
        RECT 136.600 113.800 137.000 114.200 ;
        RECT 147.800 116.200 148.200 116.600 ;
        RECT 149.400 115.500 149.800 115.900 ;
        RECT 149.400 113.100 149.800 113.500 ;
        RECT 160.600 117.800 161.000 118.200 ;
        RECT 155.000 114.800 155.400 115.200 ;
        RECT 152.600 113.800 153.000 114.200 ;
        RECT 151.000 112.800 151.400 113.200 ;
        RECT 151.800 113.100 152.200 113.500 ;
        RECT 150.200 111.800 150.600 112.200 ;
        RECT 161.400 114.800 161.800 115.200 ;
        RECT 162.200 114.800 162.600 115.200 ;
        RECT 171.000 114.800 171.400 115.200 ;
        RECT 0.600 105.100 1.000 105.500 ;
        RECT 11.000 106.800 11.400 107.200 ;
        RECT 16.600 106.800 17.000 107.200 ;
        RECT 38.200 108.800 38.600 109.200 ;
        RECT 13.400 105.800 13.800 106.200 ;
        RECT 18.200 105.900 18.600 106.300 ;
        RECT 15.800 105.100 16.200 105.500 ;
        RECT 9.400 101.800 9.800 102.200 ;
        RECT 26.200 106.800 26.600 107.200 ;
        RECT 30.200 106.800 30.600 107.200 ;
        RECT 28.600 105.800 29.000 106.200 ;
        RECT 29.400 105.100 29.800 105.500 ;
        RECT 27.800 102.800 28.200 103.200 ;
        RECT 51.000 108.800 51.400 109.200 ;
        RECT 54.200 108.800 54.600 109.200 ;
        RECT 43.000 104.800 43.400 105.200 ;
        RECT 59.800 108.800 60.200 109.200 ;
        RECT 55.000 106.800 55.400 107.200 ;
        RECT 52.600 105.800 53.000 106.200 ;
        RECT 48.600 104.800 49.000 105.200 ;
        RECT 55.800 105.800 56.200 106.200 ;
        RECT 56.600 105.800 57.000 106.200 ;
        RECT 60.600 106.800 61.000 107.200 ;
        RECT 67.800 108.800 68.200 109.200 ;
        RECT 61.400 105.800 61.800 106.200 ;
        RECT 65.400 104.800 65.800 105.200 ;
        RECT 63.000 101.800 63.400 102.200 ;
        RECT 75.800 106.800 76.200 107.200 ;
        RECT 85.400 108.800 85.800 109.200 ;
        RECT 70.200 106.100 70.600 106.500 ;
        RECT 76.600 105.100 77.000 105.500 ;
        RECT 87.000 105.800 87.400 106.200 ;
        RECT 87.800 104.800 88.200 105.200 ;
        RECT 103.800 108.800 104.200 109.200 ;
        RECT 91.000 106.800 91.400 107.200 ;
        RECT 99.800 106.800 100.200 107.200 ;
        RECT 102.200 105.800 102.600 106.200 ;
        RECT 92.600 101.800 93.000 102.200 ;
        RECT 107.000 108.800 107.400 109.200 ;
        RECT 106.200 106.800 106.600 107.200 ;
        RECT 109.400 105.800 109.800 106.200 ;
        RECT 103.800 101.800 104.200 102.200 ;
        RECT 110.200 101.800 110.600 102.200 ;
        RECT 111.000 108.800 111.400 109.200 ;
        RECT 121.400 106.800 121.800 107.200 ;
        RECT 113.400 106.100 113.800 106.500 ;
        RECT 123.000 105.900 123.400 106.300 ;
        RECT 119.800 105.100 120.200 105.500 ;
        RECT 120.600 105.100 121.000 105.500 ;
        RECT 131.000 106.800 131.400 107.200 ;
        RECT 135.800 106.800 136.200 107.200 ;
        RECT 134.200 105.800 134.600 106.200 ;
        RECT 129.400 101.800 129.800 102.200 ;
        RECT 130.200 105.100 130.600 105.500 ;
        RECT 143.800 105.800 144.200 106.200 ;
        RECT 161.400 108.800 161.800 109.200 ;
        RECT 164.600 108.800 165.000 109.200 ;
        RECT 167.800 108.800 168.200 109.200 ;
        RECT 165.400 106.800 165.800 107.200 ;
        RECT 151.800 106.100 152.200 106.500 ;
        RECT 155.800 105.900 156.200 106.300 ;
        RECT 158.200 105.100 158.600 105.500 ;
        RECT 149.400 103.800 149.800 104.200 ;
        RECT 161.400 104.800 161.800 105.200 ;
        RECT 167.000 106.800 167.400 107.200 ;
        RECT 170.200 105.800 170.600 106.200 ;
        RECT 176.600 106.800 177.000 107.200 ;
        RECT 173.400 106.100 173.800 106.500 ;
        RECT 179.800 105.100 180.200 105.500 ;
        RECT 9.400 96.800 9.800 97.200 ;
        RECT 3.800 94.800 4.200 95.200 ;
        RECT 0.600 93.100 1.000 93.500 ;
        RECT 3.000 92.800 3.400 93.200 ;
        RECT 15.000 94.800 15.400 95.200 ;
        RECT 15.800 94.800 16.200 95.200 ;
        RECT 20.600 93.800 21.000 94.200 ;
        RECT 19.000 91.800 19.400 92.200 ;
        RECT 22.200 92.800 22.600 93.200 ;
        RECT 33.400 96.200 33.800 96.600 ;
        RECT 37.400 96.800 37.800 97.200 ;
        RECT 35.000 95.500 35.400 95.900 ;
        RECT 35.800 95.800 36.200 96.200 ;
        RECT 45.400 98.800 45.800 99.200 ;
        RECT 47.800 98.800 48.200 99.200 ;
        RECT 51.000 98.800 51.400 99.200 ;
        RECT 44.600 96.800 45.000 97.200 ;
        RECT 48.600 96.800 49.000 97.200 ;
        RECT 35.000 93.100 35.400 93.500 ;
        RECT 26.200 91.800 26.600 92.200 ;
        RECT 46.200 95.800 46.600 96.200 ;
        RECT 47.000 95.800 47.400 96.200 ;
        RECT 45.400 94.800 45.800 95.200 ;
        RECT 43.000 91.800 43.400 92.200 ;
        RECT 51.800 93.800 52.200 94.200 ;
        RECT 67.800 98.800 68.200 99.200 ;
        RECT 57.400 94.800 57.800 95.200 ;
        RECT 62.200 94.800 62.600 95.200 ;
        RECT 56.600 93.800 57.000 94.200 ;
        RECT 59.800 93.800 60.200 94.200 ;
        RECT 57.400 92.800 57.800 93.200 ;
        RECT 59.000 93.100 59.400 93.500 ;
        RECT 56.600 91.800 57.000 92.200 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 82.200 96.200 82.600 96.600 ;
        RECT 83.800 95.500 84.200 95.900 ;
        RECT 86.200 98.800 86.600 99.200 ;
        RECT 93.400 96.200 93.800 96.600 ;
        RECT 95.000 95.500 95.400 95.900 ;
        RECT 96.600 98.800 97.000 99.200 ;
        RECT 95.800 93.800 96.200 94.200 ;
        RECT 83.800 93.100 84.200 93.500 ;
        RECT 75.000 91.800 75.400 92.200 ;
        RECT 95.000 93.100 95.400 93.500 ;
        RECT 98.200 93.800 98.600 94.200 ;
        RECT 100.600 98.800 101.000 99.200 ;
        RECT 107.800 96.200 108.200 96.600 ;
        RECT 112.600 98.800 113.000 99.200 ;
        RECT 109.400 95.500 109.800 95.900 ;
        RECT 99.800 91.800 100.200 92.200 ;
        RECT 113.400 94.800 113.800 95.200 ;
        RECT 114.200 94.800 114.600 95.200 ;
        RECT 123.800 97.200 124.200 97.600 ;
        RECT 125.400 97.500 125.800 97.900 ;
        RECT 123.000 96.200 123.400 96.600 ;
        RECT 109.400 93.100 109.800 93.500 ;
        RECT 118.200 92.800 118.600 93.200 ;
        RECT 127.800 93.800 128.200 94.200 ;
        RECT 126.200 92.800 126.600 93.200 ;
        RECT 123.000 92.100 123.400 92.500 ;
        RECT 123.800 92.100 124.200 92.500 ;
        RECT 124.600 92.100 125.000 92.500 ;
        RECT 125.400 92.100 125.800 92.500 ;
        RECT 127.000 92.100 127.400 92.500 ;
        RECT 128.600 92.100 129.000 92.500 ;
        RECT 129.400 92.100 129.800 92.500 ;
        RECT 130.200 92.100 130.600 92.500 ;
        RECT 145.400 97.500 145.800 97.900 ;
        RECT 143.800 96.800 144.200 97.200 ;
        RECT 146.200 96.200 146.600 96.600 ;
        RECT 140.600 94.100 141.000 94.500 ;
        RECT 145.400 94.300 145.800 94.700 ;
        RECT 143.000 93.800 143.400 94.200 ;
        RECT 140.600 92.100 141.000 92.500 ;
        RECT 141.400 92.100 141.800 92.500 ;
        RECT 142.200 92.100 142.600 92.500 ;
        RECT 143.800 92.100 144.200 92.500 ;
        RECT 145.400 92.100 145.800 92.500 ;
        RECT 146.200 92.100 146.600 92.500 ;
        RECT 147.000 92.100 147.400 92.500 ;
        RECT 147.800 92.100 148.200 92.500 ;
        RECT 160.600 95.800 161.000 96.200 ;
        RECT 157.400 94.800 157.800 95.200 ;
        RECT 158.200 94.800 158.600 95.200 ;
        RECT 162.200 94.800 162.600 95.200 ;
        RECT 163.000 94.800 163.400 95.200 ;
        RECT 164.600 94.800 165.000 95.200 ;
        RECT 152.600 91.800 153.000 92.200 ;
        RECT 172.600 96.200 173.000 96.600 ;
        RECT 174.200 95.500 174.600 95.900 ;
        RECT 175.000 94.800 175.400 95.200 ;
        RECT 177.400 94.800 177.800 95.200 ;
        RECT 174.200 93.100 174.600 93.500 ;
        RECT 9.400 88.800 9.800 89.200 ;
        RECT 0.600 85.100 1.000 85.500 ;
        RECT 12.600 85.800 13.000 86.200 ;
        RECT 17.400 84.800 17.800 85.200 ;
        RECT 20.600 86.800 21.000 87.200 ;
        RECT 18.200 81.800 18.600 82.200 ;
        RECT 25.400 85.800 25.800 86.200 ;
        RECT 23.000 84.800 23.400 85.200 ;
        RECT 27.000 84.800 27.400 85.200 ;
        RECT 22.200 81.800 22.600 82.200 ;
        RECT 29.400 86.800 29.800 87.200 ;
        RECT 42.200 88.800 42.600 89.200 ;
        RECT 47.000 88.800 47.400 89.200 ;
        RECT 37.400 85.800 37.800 86.200 ;
        RECT 35.000 84.800 35.400 85.200 ;
        RECT 43.000 86.800 43.400 87.200 ;
        RECT 40.600 85.800 41.000 86.200 ;
        RECT 43.800 85.800 44.200 86.200 ;
        RECT 27.800 81.800 28.200 82.200 ;
        RECT 39.000 81.800 39.400 82.200 ;
        RECT 58.200 88.800 58.600 89.200 ;
        RECT 55.000 86.800 55.400 87.200 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 49.400 86.100 49.800 86.500 ;
        RECT 46.200 84.800 46.600 85.200 ;
        RECT 53.400 85.900 53.800 86.300 ;
        RECT 55.800 85.100 56.200 85.500 ;
        RECT 61.400 85.800 61.800 86.200 ;
        RECT 73.400 88.800 73.800 89.200 ;
        RECT 66.200 85.800 66.600 86.200 ;
        RECT 63.800 84.800 64.200 85.200 ;
        RECT 63.000 81.800 63.400 82.200 ;
        RECT 69.400 84.800 69.800 85.200 ;
        RECT 71.800 85.800 72.200 86.200 ;
        RECT 84.600 88.800 85.000 89.200 ;
        RECT 74.200 86.800 74.600 87.200 ;
        RECT 75.000 85.800 75.400 86.200 ;
        RECT 79.000 85.800 79.400 86.200 ;
        RECT 80.600 84.800 81.000 85.200 ;
        RECT 78.200 81.800 78.600 82.200 ;
        RECT 91.000 88.800 91.400 89.200 ;
        RECT 96.600 88.800 97.000 89.200 ;
        RECT 84.600 84.800 85.000 85.200 ;
        RECT 93.400 85.800 93.800 86.200 ;
        RECT 95.000 85.800 95.400 86.200 ;
        RECT 101.400 87.800 101.800 88.200 ;
        RECT 99.000 86.800 99.400 87.200 ;
        RECT 98.200 85.800 98.600 86.200 ;
        RECT 99.800 85.800 100.200 86.200 ;
        RECT 106.200 85.900 106.600 86.300 ;
        RECT 103.800 85.100 104.200 85.500 ;
        RECT 115.800 88.800 116.200 89.200 ;
        RECT 120.600 88.800 121.000 89.200 ;
        RECT 116.600 86.800 117.000 87.200 ;
        RECT 117.400 85.800 117.800 86.200 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 114.200 81.800 114.600 82.200 ;
        RECT 123.800 84.800 124.200 85.200 ;
        RECT 124.600 85.100 125.000 85.500 ;
        RECT 135.800 88.800 136.200 89.200 ;
        RECT 135.000 86.800 135.400 87.200 ;
        RECT 140.600 87.800 141.000 88.200 ;
        RECT 137.400 85.800 137.800 86.200 ;
        RECT 145.400 86.500 145.800 86.900 ;
        RECT 133.400 81.800 133.800 82.200 ;
        RECT 150.200 86.300 150.600 86.700 ;
        RECT 157.400 87.800 157.800 88.200 ;
        RECT 160.600 88.800 161.000 89.200 ;
        RECT 159.800 86.800 160.200 87.200 ;
        RECT 167.800 86.800 168.200 87.200 ;
        RECT 173.400 87.800 173.800 88.200 ;
        RECT 162.200 85.800 162.600 86.200 ;
        RECT 146.200 84.400 146.600 84.800 ;
        RECT 148.600 83.800 149.000 84.200 ;
        RECT 147.000 83.100 147.400 83.500 ;
        RECT 145.400 82.100 145.800 82.500 ;
        RECT 146.200 82.100 146.600 82.500 ;
        RECT 148.600 83.100 149.000 83.500 ;
        RECT 150.200 83.100 150.600 83.500 ;
        RECT 151.000 82.100 151.400 82.500 ;
        RECT 151.800 82.100 152.200 82.500 ;
        RECT 152.600 82.100 153.000 82.500 ;
        RECT 171.000 84.800 171.400 85.200 ;
        RECT 3.800 74.800 4.200 75.200 ;
        RECT 0.600 73.100 1.000 73.500 ;
        RECT 9.400 71.800 9.800 72.200 ;
        RECT 12.600 76.800 13.000 77.200 ;
        RECT 11.000 72.800 11.400 73.200 ;
        RECT 10.200 71.800 10.600 72.200 ;
        RECT 14.200 72.800 14.600 73.200 ;
        RECT 21.400 78.800 21.800 79.200 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 19.800 74.800 20.200 75.200 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 25.400 78.800 25.800 79.200 ;
        RECT 23.000 76.800 23.400 77.200 ;
        RECT 24.600 76.800 25.000 77.200 ;
        RECT 23.000 75.800 23.400 76.200 ;
        RECT 35.000 78.800 35.400 79.200 ;
        RECT 29.400 74.800 29.800 75.200 ;
        RECT 26.200 73.100 26.600 73.500 ;
        RECT 44.600 78.800 45.000 79.200 ;
        RECT 42.200 74.800 42.600 75.200 ;
        RECT 43.000 74.800 43.400 75.200 ;
        RECT 43.800 73.800 44.200 74.200 ;
        RECT 49.400 74.800 49.800 75.200 ;
        RECT 47.000 73.800 47.400 74.200 ;
        RECT 46.200 73.100 46.600 73.500 ;
        RECT 57.400 73.800 57.800 74.200 ;
        RECT 65.400 76.200 65.800 76.600 ;
        RECT 67.000 75.500 67.400 75.900 ;
        RECT 74.200 78.800 74.600 79.200 ;
        RECT 55.000 71.800 55.400 72.200 ;
        RECT 64.600 72.800 65.000 73.200 ;
        RECT 67.000 73.100 67.400 73.500 ;
        RECT 67.800 72.800 68.200 73.200 ;
        RECT 76.600 76.800 77.000 77.200 ;
        RECT 72.600 74.800 73.000 75.200 ;
        RECT 73.400 74.800 73.800 75.200 ;
        RECT 75.800 74.800 76.200 75.200 ;
        RECT 79.000 78.800 79.400 79.200 ;
        RECT 78.200 73.800 78.600 74.200 ;
        RECT 81.400 73.800 81.800 74.200 ;
        RECT 93.400 76.200 93.800 76.600 ;
        RECT 95.000 75.500 95.400 75.900 ;
        RECT 96.600 78.800 97.000 79.200 ;
        RECT 95.800 73.800 96.200 74.200 ;
        RECT 95.000 73.100 95.400 73.500 ;
        RECT 86.200 71.800 86.600 72.200 ;
        RECT 105.400 74.800 105.800 75.200 ;
        RECT 106.200 74.800 106.600 75.200 ;
        RECT 97.400 71.800 97.800 72.200 ;
        RECT 100.600 73.800 101.000 74.200 ;
        RECT 113.400 77.800 113.800 78.200 ;
        RECT 111.000 74.800 111.400 75.200 ;
        RECT 103.000 72.800 103.400 73.200 ;
        RECT 104.600 72.800 105.000 73.200 ;
        RECT 101.400 71.800 101.800 72.200 ;
        RECT 112.600 73.800 113.000 74.200 ;
        RECT 107.800 71.800 108.200 72.200 ;
        RECT 115.800 78.800 116.200 79.200 ;
        RECT 123.000 76.800 123.400 77.200 ;
        RECT 115.800 73.800 116.200 74.200 ;
        RECT 115.800 72.800 116.200 73.200 ;
        RECT 118.200 74.800 118.600 75.200 ;
        RECT 122.200 74.800 122.600 75.200 ;
        RECT 123.800 74.800 124.200 75.200 ;
        RECT 125.400 74.800 125.800 75.200 ;
        RECT 126.200 74.800 126.600 75.200 ;
        RECT 124.600 73.800 125.000 74.200 ;
        RECT 129.400 73.800 129.800 74.200 ;
        RECT 138.200 76.800 138.600 77.200 ;
        RECT 135.000 74.800 135.400 75.200 ;
        RECT 137.400 74.800 137.800 75.200 ;
        RECT 131.000 72.800 131.400 73.200 ;
        RECT 145.400 76.200 145.800 76.600 ;
        RECT 147.000 75.500 147.400 75.900 ;
        RECT 156.600 77.500 157.000 77.900 ;
        RECT 155.000 76.800 155.400 77.200 ;
        RECT 157.400 76.200 157.800 76.600 ;
        RECT 151.800 74.100 152.200 74.500 ;
        RECT 156.600 74.300 157.000 74.700 ;
        RECT 144.600 72.800 145.000 73.200 ;
        RECT 147.000 73.100 147.400 73.500 ;
        RECT 154.200 73.800 154.600 74.200 ;
        RECT 151.800 72.100 152.200 72.500 ;
        RECT 152.600 72.100 153.000 72.500 ;
        RECT 153.400 72.100 153.800 72.500 ;
        RECT 155.000 72.100 155.400 72.500 ;
        RECT 156.600 72.100 157.000 72.500 ;
        RECT 157.400 72.100 157.800 72.500 ;
        RECT 158.200 72.100 158.600 72.500 ;
        RECT 159.000 72.100 159.400 72.500 ;
        RECT 170.200 78.800 170.600 79.200 ;
        RECT 165.400 74.800 165.800 75.200 ;
        RECT 166.200 74.800 166.600 75.200 ;
        RECT 169.400 74.800 169.800 75.200 ;
        RECT 168.600 73.800 169.000 74.200 ;
        RECT 163.800 71.800 164.200 72.200 ;
        RECT 177.400 76.200 177.800 76.600 ;
        RECT 179.000 75.500 179.400 75.900 ;
        RECT 179.000 73.100 179.400 73.500 ;
        RECT 9.400 68.800 9.800 69.200 ;
        RECT 7.800 66.800 8.200 67.200 ;
        RECT 3.000 61.800 3.400 62.200 ;
        RECT 8.600 65.800 9.000 66.200 ;
        RECT 15.800 66.800 16.200 67.200 ;
        RECT 11.800 66.100 12.200 66.500 ;
        RECT 23.800 66.800 24.200 67.200 ;
        RECT 18.200 65.100 18.600 65.500 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 23.800 64.800 24.200 65.200 ;
        RECT 27.800 68.800 28.200 69.200 ;
        RECT 27.000 66.800 27.400 67.200 ;
        RECT 39.000 68.800 39.400 69.200 ;
        RECT 38.200 66.800 38.600 67.200 ;
        RECT 30.200 66.100 30.600 66.500 ;
        RECT 31.800 65.800 32.200 66.200 ;
        RECT 47.000 66.800 47.400 67.200 ;
        RECT 41.400 66.100 41.800 66.500 ;
        RECT 45.400 65.900 45.800 66.300 ;
        RECT 36.600 65.100 37.000 65.500 ;
        RECT 47.800 65.100 48.200 65.500 ;
        RECT 53.400 65.800 53.800 66.200 ;
        RECT 63.800 68.800 64.200 69.200 ;
        RECT 62.200 65.800 62.600 66.200 ;
        RECT 67.000 68.800 67.400 69.200 ;
        RECT 64.600 66.800 65.000 67.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 69.400 68.800 69.800 69.200 ;
        RECT 79.000 68.800 79.400 69.200 ;
        RECT 70.200 65.100 70.600 65.500 ;
        RECT 91.000 66.800 91.400 67.200 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 89.400 65.800 89.800 66.200 ;
        RECT 94.200 66.100 94.600 66.500 ;
        RECT 98.200 65.900 98.600 66.300 ;
        RECT 116.600 68.800 117.000 69.200 ;
        RECT 100.600 65.100 101.000 65.500 ;
        RECT 107.800 65.100 108.200 65.500 ;
        RECT 119.000 65.800 119.400 66.200 ;
        RECT 123.000 66.800 123.400 67.200 ;
        RECT 123.800 65.800 124.200 66.200 ;
        RECT 127.000 65.900 127.400 66.300 ;
        RECT 124.600 65.100 125.000 65.500 ;
        RECT 135.800 66.800 136.200 67.200 ;
        RECT 141.400 66.800 141.800 67.200 ;
        RECT 147.800 66.800 148.200 67.200 ;
        RECT 153.400 68.800 153.800 69.200 ;
        RECT 151.800 66.800 152.200 67.200 ;
        RECT 152.600 66.800 153.000 67.200 ;
        RECT 143.800 64.800 144.200 65.200 ;
        RECT 158.200 65.800 158.600 66.200 ;
        RECT 163.000 66.800 163.400 67.200 ;
        RECT 179.800 68.800 180.200 69.200 ;
        RECT 167.000 65.800 167.400 66.200 ;
        RECT 174.200 66.800 174.600 67.200 ;
        RECT 171.800 66.100 172.200 66.500 ;
        RECT 178.200 65.100 178.600 65.500 ;
        RECT 169.400 61.800 169.800 62.200 ;
        RECT 179.800 61.800 180.200 62.200 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 4.600 54.800 5.000 55.200 ;
        RECT 6.200 54.800 6.600 55.200 ;
        RECT 21.400 58.800 21.800 59.200 ;
        RECT 3.000 51.800 3.400 52.200 ;
        RECT 7.800 53.800 8.200 54.200 ;
        RECT 11.000 53.100 11.400 53.500 ;
        RECT 8.600 51.800 9.000 52.200 ;
        RECT 40.600 56.800 41.000 57.200 ;
        RECT 44.600 56.800 45.000 57.200 ;
        RECT 47.800 58.800 48.200 59.200 ;
        RECT 47.000 56.800 47.400 57.200 ;
        RECT 31.800 53.800 32.200 54.200 ;
        RECT 19.800 51.800 20.200 52.200 ;
        RECT 30.200 52.800 30.600 53.200 ;
        RECT 31.000 53.100 31.400 53.500 ;
        RECT 36.600 53.800 37.000 54.200 ;
        RECT 48.600 55.800 49.000 56.200 ;
        RECT 47.800 54.800 48.200 55.200 ;
        RECT 52.600 58.800 53.000 59.200 ;
        RECT 51.800 53.800 52.200 54.200 ;
        RECT 56.600 56.800 57.000 57.200 ;
        RECT 53.400 53.800 53.800 54.200 ;
        RECT 54.200 52.800 54.600 53.200 ;
        RECT 55.000 51.800 55.400 52.200 ;
        RECT 63.800 56.200 64.200 56.600 ;
        RECT 71.800 58.800 72.200 59.200 ;
        RECT 65.400 55.500 65.800 55.900 ;
        RECT 65.400 53.100 65.800 53.500 ;
        RECT 67.800 52.800 68.200 53.200 ;
        RECT 68.600 52.800 69.000 53.200 ;
        RECT 73.400 54.800 73.800 55.200 ;
        RECT 74.200 54.800 74.600 55.200 ;
        RECT 82.200 58.800 82.600 59.200 ;
        RECT 83.800 58.800 84.200 59.200 ;
        RECT 72.600 52.800 73.000 53.200 ;
        RECT 79.800 53.800 80.200 54.200 ;
        RECT 91.000 56.200 91.400 56.600 ;
        RECT 100.600 58.800 101.000 59.200 ;
        RECT 92.600 55.500 93.000 55.900 ;
        RECT 92.600 53.100 93.000 53.500 ;
        RECT 96.600 52.800 97.000 53.200 ;
        RECT 98.200 52.800 98.600 53.200 ;
        RECT 107.800 56.200 108.200 56.600 ;
        RECT 109.400 55.500 109.800 55.900 ;
        RECT 109.400 53.100 109.800 53.500 ;
        RECT 110.200 52.800 110.600 53.200 ;
        RECT 117.400 58.800 117.800 59.200 ;
        RECT 115.000 54.800 115.400 55.200 ;
        RECT 115.800 54.800 116.200 55.200 ;
        RECT 116.600 52.800 117.000 53.200 ;
        RECT 119.000 58.800 119.400 59.200 ;
        RECT 118.200 53.800 118.600 54.200 ;
        RECT 121.400 58.800 121.800 59.200 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 124.600 53.800 125.000 54.200 ;
        RECT 134.200 56.200 134.600 56.600 ;
        RECT 135.800 55.500 136.200 55.900 ;
        RECT 138.200 55.800 138.600 56.200 ;
        RECT 126.200 52.800 126.600 53.200 ;
        RECT 135.800 53.100 136.200 53.500 ;
        RECT 127.000 51.800 127.400 52.200 ;
        RECT 136.600 52.800 137.000 53.200 ;
        RECT 143.000 54.800 143.400 55.200 ;
        RECT 143.800 54.800 144.200 55.200 ;
        RECT 147.800 54.800 148.200 55.200 ;
        RECT 167.800 58.800 168.200 59.200 ;
        RECT 170.200 58.800 170.600 59.200 ;
        RECT 145.400 53.800 145.800 54.200 ;
        RECT 144.600 53.100 145.000 53.500 ;
        RECT 150.200 53.800 150.600 54.200 ;
        RECT 154.200 54.800 154.600 55.200 ;
        RECT 155.000 54.800 155.400 55.200 ;
        RECT 163.000 55.700 163.400 56.100 ;
        RECT 153.400 51.800 153.800 52.200 ;
        RECT 165.400 54.800 165.800 55.200 ;
        RECT 166.200 54.800 166.600 55.200 ;
        RECT 156.600 51.800 157.000 52.200 ;
        RECT 177.400 56.200 177.800 56.600 ;
        RECT 179.000 55.500 179.400 55.900 ;
        RECT 174.200 54.800 174.600 55.200 ;
        RECT 179.000 53.100 179.400 53.500 ;
        RECT 9.400 48.800 9.800 49.200 ;
        RECT 3.000 45.900 3.400 46.300 ;
        RECT 0.600 45.100 1.000 45.500 ;
        RECT 21.400 48.800 21.800 49.200 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 11.000 41.800 11.400 42.200 ;
        RECT 31.800 46.800 32.200 47.200 ;
        RECT 19.800 44.800 20.200 45.200 ;
        RECT 35.000 47.800 35.400 48.200 ;
        RECT 44.600 48.800 45.000 49.200 ;
        RECT 36.600 46.800 37.000 47.200 ;
        RECT 38.200 45.900 38.600 46.300 ;
        RECT 35.800 45.100 36.200 45.500 ;
        RECT 51.000 48.800 51.400 49.200 ;
        RECT 55.800 48.800 56.200 49.200 ;
        RECT 54.200 45.800 54.600 46.200 ;
        RECT 64.600 48.800 65.000 49.200 ;
        RECT 68.600 48.800 69.000 49.200 ;
        RECT 58.200 46.800 58.600 47.200 ;
        RECT 60.600 46.800 61.000 47.200 ;
        RECT 57.400 45.800 57.800 46.200 ;
        RECT 58.200 45.800 58.600 46.200 ;
        RECT 64.600 46.800 65.000 47.200 ;
        RECT 63.800 45.800 64.200 46.200 ;
        RECT 66.200 45.800 66.600 46.200 ;
        RECT 79.800 48.800 80.200 49.200 ;
        RECT 71.800 46.800 72.200 47.200 ;
        RECT 90.200 48.800 90.600 49.200 ;
        RECT 75.000 45.800 75.400 46.200 ;
        RECT 71.000 45.100 71.400 45.500 ;
        RECT 81.400 46.800 81.800 47.200 ;
        RECT 80.600 45.100 81.000 45.500 ;
        RECT 87.800 43.800 88.200 44.200 ;
        RECT 100.600 48.800 101.000 49.200 ;
        RECT 103.800 48.800 104.200 49.200 ;
        RECT 99.000 46.800 99.400 47.200 ;
        RECT 101.400 45.800 101.800 46.200 ;
        RECT 105.400 45.800 105.800 46.200 ;
        RECT 108.600 48.800 109.000 49.200 ;
        RECT 107.000 41.800 107.400 42.200 ;
        RECT 118.200 48.800 118.600 49.200 ;
        RECT 110.200 46.800 110.600 47.200 ;
        RECT 119.000 48.800 119.400 49.200 ;
        RECT 109.400 45.100 109.800 45.500 ;
        RECT 126.200 48.800 126.600 49.200 ;
        RECT 132.600 48.800 133.000 49.200 ;
        RECT 124.600 45.800 125.000 46.200 ;
        RECT 127.800 45.800 128.200 46.200 ;
        RECT 126.200 44.800 126.600 45.200 ;
        RECT 142.200 48.800 142.600 49.200 ;
        RECT 140.600 47.800 141.000 48.200 ;
        RECT 135.800 41.800 136.200 42.200 ;
        RECT 155.800 48.800 156.200 49.200 ;
        RECT 156.600 48.800 157.000 49.200 ;
        RECT 151.800 45.800 152.200 46.200 ;
        RECT 168.600 48.800 169.000 49.200 ;
        RECT 169.400 48.800 169.800 49.200 ;
        RECT 159.000 46.100 159.400 46.500 ;
        RECT 151.000 41.800 151.400 42.200 ;
        RECT 155.800 44.800 156.200 45.200 ;
        RECT 165.400 45.100 165.800 45.500 ;
        RECT 168.600 44.800 169.000 45.200 ;
        RECT 173.400 46.100 173.800 46.500 ;
        RECT 179.800 45.100 180.200 45.500 ;
        RECT 171.000 41.800 171.400 42.200 ;
        RECT 9.400 38.800 9.800 39.200 ;
        RECT 3.800 34.800 4.200 35.200 ;
        RECT 0.600 33.100 1.000 33.500 ;
        RECT 17.400 38.800 17.800 39.200 ;
        RECT 27.800 36.800 28.200 37.200 ;
        RECT 13.400 34.800 13.800 35.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 22.200 34.800 22.600 35.200 ;
        RECT 3.000 32.800 3.400 33.200 ;
        RECT 19.000 33.100 19.400 33.500 ;
        RECT 28.600 34.800 29.000 35.200 ;
        RECT 29.400 34.800 29.800 35.200 ;
        RECT 21.400 32.800 21.800 33.200 ;
        RECT 35.000 34.800 35.400 35.200 ;
        RECT 35.800 34.800 36.200 35.200 ;
        RECT 44.600 38.800 45.000 39.200 ;
        RECT 50.200 38.800 50.600 39.200 ;
        RECT 43.800 36.800 44.200 37.200 ;
        RECT 47.800 36.800 48.200 37.200 ;
        RECT 34.200 32.800 34.600 33.200 ;
        RECT 37.400 31.800 37.800 32.200 ;
        RECT 51.000 36.800 51.400 37.200 ;
        RECT 46.200 35.800 46.600 36.200 ;
        RECT 44.600 34.800 45.000 35.200 ;
        RECT 42.200 32.800 42.600 33.200 ;
        RECT 55.000 38.800 55.400 39.200 ;
        RECT 55.800 36.800 56.200 37.200 ;
        RECT 54.200 35.800 54.600 36.200 ;
        RECT 65.400 38.800 65.800 39.200 ;
        RECT 59.000 34.800 59.400 35.200 ;
        RECT 52.600 33.800 53.000 34.200 ;
        RECT 53.400 33.800 53.800 34.200 ;
        RECT 59.000 32.800 59.400 33.200 ;
        RECT 71.800 38.800 72.200 39.200 ;
        RECT 81.400 38.800 81.800 39.200 ;
        RECT 79.800 37.800 80.200 38.200 ;
        RECT 83.800 36.800 84.200 37.200 ;
        RECT 79.000 31.800 79.400 32.200 ;
        RECT 87.000 34.800 87.400 35.200 ;
        RECT 88.600 34.800 89.000 35.200 ;
        RECT 82.200 32.800 82.600 33.200 ;
        RECT 89.400 34.800 89.800 35.200 ;
        RECT 103.800 38.800 104.200 39.200 ;
        RECT 110.200 36.800 110.600 37.200 ;
        RECT 95.800 33.800 96.200 34.200 ;
        RECT 94.200 32.800 94.600 33.200 ;
        RECT 95.000 33.100 95.400 33.500 ;
        RECT 104.600 32.800 105.000 33.200 ;
        RECT 107.800 32.800 108.200 33.200 ;
        RECT 117.400 36.200 117.800 36.600 ;
        RECT 119.000 35.500 119.400 35.900 ;
        RECT 120.600 34.800 121.000 35.200 ;
        RECT 125.400 38.800 125.800 39.200 ;
        RECT 119.000 33.100 119.400 33.500 ;
        RECT 123.000 32.800 123.400 33.200 ;
        RECT 142.200 38.800 142.600 39.200 ;
        RECT 146.200 38.800 146.600 39.200 ;
        RECT 134.200 33.800 134.600 34.200 ;
        RECT 125.400 31.800 125.800 32.200 ;
        RECT 127.000 31.800 127.400 32.200 ;
        RECT 133.400 33.100 133.800 33.500 ;
        RECT 146.200 34.800 146.600 35.200 ;
        RECT 151.000 34.800 151.400 35.200 ;
        RECT 147.000 33.800 147.400 34.200 ;
        RECT 147.800 33.100 148.200 33.500 ;
        RECT 158.200 38.800 158.600 39.200 ;
        RECT 162.200 34.800 162.600 35.200 ;
        RECT 159.000 32.800 159.400 33.200 ;
        RECT 163.800 34.800 164.200 35.200 ;
        RECT 164.600 34.800 165.000 35.200 ;
        RECT 172.600 36.200 173.000 36.600 ;
        RECT 174.200 35.500 174.600 35.900 ;
        RECT 169.400 34.800 169.800 35.200 ;
        RECT 175.000 34.800 175.400 35.200 ;
        RECT 175.800 34.800 176.200 35.200 ;
        RECT 174.200 33.100 174.600 33.500 ;
        RECT 165.400 31.800 165.800 32.200 ;
        RECT 9.400 28.800 9.800 29.200 ;
        RECT 0.600 25.100 1.000 25.500 ;
        RECT 19.000 28.800 19.400 29.200 ;
        RECT 21.400 28.800 21.800 29.200 ;
        RECT 17.400 26.800 17.800 27.200 ;
        RECT 36.600 28.800 37.000 29.200 ;
        RECT 19.800 25.800 20.200 26.200 ;
        RECT 28.600 26.800 29.000 27.200 ;
        RECT 40.600 28.800 41.000 29.200 ;
        RECT 27.800 25.100 28.200 25.500 ;
        RECT 44.600 26.800 45.000 27.200 ;
        RECT 44.600 25.800 45.000 26.200 ;
        RECT 42.200 23.800 42.600 24.200 ;
        RECT 45.400 24.800 45.800 25.200 ;
        RECT 53.400 28.800 53.800 29.200 ;
        RECT 49.400 25.800 49.800 26.200 ;
        RECT 57.400 28.800 57.800 29.200 ;
        RECT 54.200 25.800 54.600 26.200 ;
        RECT 49.400 21.800 49.800 22.200 ;
        RECT 65.400 28.800 65.800 29.200 ;
        RECT 64.600 24.800 65.000 25.200 ;
        RECT 68.600 28.800 69.000 29.200 ;
        RECT 75.800 28.800 76.200 29.200 ;
        RECT 79.800 28.800 80.200 29.200 ;
        RECT 76.600 27.800 77.000 28.200 ;
        RECT 75.000 25.800 75.400 26.200 ;
        RECT 77.400 25.800 77.800 26.200 ;
        RECT 82.200 28.800 82.600 29.200 ;
        RECT 87.800 26.800 88.200 27.200 ;
        RECT 84.600 26.100 85.000 26.500 ;
        RECT 88.600 25.900 89.000 26.300 ;
        RECT 91.000 25.100 91.400 25.500 ;
        RECT 99.800 25.800 100.200 26.200 ;
        RECT 103.800 26.800 104.200 27.200 ;
        RECT 116.600 28.800 117.000 29.200 ;
        RECT 114.200 26.800 114.600 27.200 ;
        RECT 108.600 26.100 109.000 26.500 ;
        RECT 115.000 25.100 115.400 25.500 ;
        RECT 115.800 24.800 116.200 25.200 ;
        RECT 122.200 26.800 122.600 27.200 ;
        RECT 125.400 28.800 125.800 29.200 ;
        RECT 124.600 24.800 125.000 25.200 ;
        RECT 136.600 28.800 137.000 29.200 ;
        RECT 142.200 28.800 142.600 29.200 ;
        RECT 129.400 26.100 129.800 26.500 ;
        RECT 135.800 25.100 136.200 25.500 ;
        RECT 140.600 25.800 141.000 26.200 ;
        RECT 141.400 24.800 141.800 25.200 ;
        RECT 144.600 21.800 145.000 22.200 ;
        RECT 145.400 28.800 145.800 29.200 ;
        RECT 155.800 28.800 156.200 29.200 ;
        RECT 147.800 26.100 148.200 26.500 ;
        RECT 149.400 25.800 149.800 26.200 ;
        RECT 154.200 25.100 154.600 25.500 ;
        RECT 156.600 24.800 157.000 25.200 ;
        RECT 169.400 28.800 169.800 29.200 ;
        RECT 161.400 26.800 161.800 27.200 ;
        RECT 164.600 25.800 165.000 26.200 ;
        RECT 159.000 21.800 159.400 22.200 ;
        RECT 160.600 25.100 161.000 25.500 ;
        RECT 170.200 28.800 170.600 29.200 ;
        RECT 171.800 28.800 172.200 29.200 ;
        RECT 177.400 28.800 177.800 29.200 ;
        RECT 178.200 24.800 178.600 25.200 ;
        RECT 6.200 15.800 6.600 16.200 ;
        RECT 12.600 18.800 13.000 19.200 ;
        RECT 3.800 14.800 4.200 15.200 ;
        RECT 4.600 14.800 5.000 15.200 ;
        RECT 3.000 11.800 3.400 12.200 ;
        RECT 6.200 12.800 6.600 13.200 ;
        RECT 19.800 16.200 20.200 16.600 ;
        RECT 21.400 15.500 21.800 15.900 ;
        RECT 22.200 14.800 22.600 15.200 ;
        RECT 23.000 14.800 23.400 15.200 ;
        RECT 37.400 16.800 37.800 17.200 ;
        RECT 8.600 11.800 9.000 12.200 ;
        RECT 11.800 12.800 12.200 13.200 ;
        RECT 15.800 12.800 16.200 13.200 ;
        RECT 21.400 13.100 21.800 13.500 ;
        RECT 24.600 11.800 25.000 12.200 ;
        RECT 31.800 14.800 32.200 15.200 ;
        RECT 29.400 13.800 29.800 14.200 ;
        RECT 27.800 12.800 28.200 13.200 ;
        RECT 28.600 13.100 29.000 13.500 ;
        RECT 39.800 14.800 40.200 15.200 ;
        RECT 40.600 14.800 41.000 15.200 ;
        RECT 46.200 18.800 46.600 19.200 ;
        RECT 53.400 16.200 53.800 16.600 ;
        RECT 55.000 15.500 55.400 15.900 ;
        RECT 49.400 12.800 49.800 13.200 ;
        RECT 52.600 12.800 53.000 13.200 ;
        RECT 55.000 13.100 55.400 13.500 ;
        RECT 55.800 12.800 56.200 13.200 ;
        RECT 59.000 12.800 59.400 13.200 ;
        RECT 61.400 12.800 61.800 13.200 ;
        RECT 68.600 18.800 69.000 19.200 ;
        RECT 66.200 14.800 66.600 15.200 ;
        RECT 67.000 14.800 67.400 15.200 ;
        RECT 78.200 18.800 78.600 19.200 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 73.400 11.800 73.800 12.200 ;
        RECT 87.000 16.200 87.400 16.600 ;
        RECT 88.600 15.500 89.000 15.900 ;
        RECT 88.600 13.100 89.000 13.500 ;
        RECT 91.000 12.800 91.400 13.200 ;
        RECT 97.400 18.800 97.800 19.200 ;
        RECT 95.800 14.800 96.200 15.200 ;
        RECT 96.600 14.800 97.000 15.200 ;
        RECT 104.600 16.200 105.000 16.600 ;
        RECT 106.200 15.500 106.600 15.900 ;
        RECT 110.200 15.800 110.600 16.200 ;
        RECT 106.200 13.100 106.600 13.500 ;
        RECT 107.000 12.800 107.400 13.200 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 112.600 14.800 113.000 15.200 ;
        RECT 113.400 12.800 113.800 13.200 ;
        RECT 115.000 14.800 115.400 15.200 ;
        RECT 115.800 14.800 116.200 15.200 ;
        RECT 119.800 12.800 120.200 13.200 ;
        RECT 121.400 14.800 121.800 15.200 ;
        RECT 122.200 14.800 122.600 15.200 ;
        RECT 129.400 14.800 129.800 15.200 ;
        RECT 127.000 13.800 127.400 14.200 ;
        RECT 126.200 13.100 126.600 13.500 ;
        RECT 136.600 18.800 137.000 19.200 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 140.600 14.800 141.000 15.200 ;
        RECT 143.000 14.800 143.400 15.200 ;
        RECT 147.000 14.800 147.400 15.200 ;
        RECT 147.800 14.800 148.200 15.200 ;
        RECT 148.600 14.800 149.000 15.200 ;
        RECT 149.400 14.800 149.800 15.200 ;
        RECT 162.200 18.800 162.600 19.200 ;
        RECT 152.600 14.800 153.000 15.200 ;
        RECT 168.600 18.800 169.000 19.200 ;
        RECT 151.800 13.800 152.200 14.200 ;
        RECT 154.200 13.800 154.600 14.200 ;
        RECT 153.400 13.100 153.800 13.500 ;
        RECT 163.000 14.800 163.400 15.200 ;
        RECT 163.800 14.800 164.200 15.200 ;
        RECT 167.800 13.800 168.200 14.200 ;
        RECT 171.000 15.800 171.400 16.200 ;
        RECT 171.000 12.800 171.400 13.200 ;
        RECT 171.800 12.800 172.200 13.200 ;
        RECT 173.400 18.800 173.800 19.200 ;
        RECT 178.200 14.800 178.600 15.200 ;
        RECT 179.000 14.800 179.400 15.200 ;
        RECT 174.200 12.800 174.600 13.200 ;
        RECT 9.400 8.800 9.800 9.200 ;
        RECT 19.000 8.800 19.400 9.200 ;
        RECT 4.600 6.800 5.000 7.200 ;
        RECT 3.000 5.900 3.400 6.300 ;
        RECT 0.600 5.100 1.000 5.500 ;
        RECT 11.000 6.800 11.400 7.200 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 12.600 5.900 13.000 6.300 ;
        RECT 10.200 5.100 10.600 5.500 ;
        RECT 21.400 8.800 21.800 9.200 ;
        RECT 20.600 6.800 21.000 7.200 ;
        RECT 34.200 8.800 34.600 9.200 ;
        RECT 45.400 8.800 45.800 9.200 ;
        RECT 29.400 6.800 29.800 7.200 ;
        RECT 24.600 5.800 25.000 6.200 ;
        RECT 27.800 5.900 28.200 6.300 ;
        RECT 25.400 5.100 25.800 5.500 ;
        RECT 37.400 6.800 37.800 7.200 ;
        RECT 41.400 5.800 41.800 6.200 ;
        RECT 36.600 5.100 37.000 5.500 ;
        RECT 47.800 5.800 48.200 6.200 ;
        RECT 60.600 8.800 61.000 9.200 ;
        RECT 50.200 6.800 50.600 7.200 ;
        RECT 52.600 6.800 53.000 7.200 ;
        RECT 51.000 5.800 51.400 6.200 ;
        RECT 51.800 5.100 52.200 5.500 ;
        RECT 63.800 8.800 64.200 9.200 ;
        RECT 65.400 8.800 65.800 9.200 ;
        RECT 83.800 8.800 84.200 9.200 ;
        RECT 78.200 6.800 78.600 7.200 ;
        RECT 67.800 6.100 68.200 6.500 ;
        RECT 71.800 5.900 72.200 6.300 ;
        RECT 74.200 5.100 74.600 5.500 ;
        RECT 75.000 5.100 75.400 5.500 ;
        RECT 95.000 8.800 95.400 9.200 ;
        RECT 96.600 8.800 97.000 9.200 ;
        RECT 107.000 8.800 107.400 9.200 ;
        RECT 104.600 6.800 105.000 7.200 ;
        RECT 99.000 6.100 99.400 6.500 ;
        RECT 103.000 5.900 103.400 6.300 ;
        RECT 105.400 5.100 105.800 5.500 ;
        RECT 117.400 8.800 117.800 9.200 ;
        RECT 111.800 6.800 112.200 7.200 ;
        RECT 112.600 5.800 113.000 6.200 ;
        RECT 108.600 5.100 109.000 5.500 ;
        RECT 121.400 5.800 121.800 6.200 ;
        RECT 127.000 6.800 127.400 7.200 ;
        RECT 126.200 5.100 126.600 5.500 ;
        RECT 135.800 6.800 136.200 7.200 ;
        RECT 159.800 8.800 160.200 9.200 ;
        RECT 137.400 4.800 137.800 5.200 ;
        RECT 146.200 5.800 146.600 6.200 ;
        RECT 150.200 6.800 150.600 7.200 ;
        RECT 169.400 8.800 169.800 9.200 ;
        RECT 154.200 6.800 154.600 7.200 ;
        RECT 149.400 5.800 149.800 6.200 ;
        RECT 153.400 5.900 153.800 6.300 ;
        RECT 151.000 5.100 151.400 5.500 ;
        RECT 161.400 6.800 161.800 7.200 ;
        RECT 179.000 8.800 179.400 9.200 ;
        RECT 160.600 5.100 161.000 5.500 ;
        RECT 171.000 6.800 171.400 7.200 ;
        RECT 172.600 5.900 173.000 6.300 ;
        RECT 170.200 5.100 170.600 5.500 ;
      LAYER metal2 ;
        RECT 1.400 168.800 1.800 169.200 ;
        RECT 15.000 169.100 15.400 169.200 ;
        RECT 15.800 169.100 16.200 169.200 ;
        RECT 1.400 168.200 1.700 168.800 ;
        RECT 1.400 167.800 1.800 168.200 ;
        RECT 6.200 166.800 6.600 167.200 ;
        RECT 6.200 166.200 6.500 166.800 ;
        RECT 3.800 165.800 4.200 166.200 ;
        RECT 5.400 165.800 5.800 166.200 ;
        RECT 6.200 165.800 6.600 166.200 ;
        RECT 3.800 165.200 4.100 165.800 ;
        RECT 3.800 164.800 4.200 165.200 ;
        RECT 0.600 153.100 1.000 155.900 ;
        RECT 2.200 152.100 2.600 157.900 ;
        RECT 5.400 155.200 5.700 165.800 ;
        RECT 7.000 165.100 7.400 167.900 ;
        RECT 8.600 163.100 9.000 168.900 ;
        RECT 9.400 165.900 9.800 166.300 ;
        RECT 9.400 165.200 9.700 165.900 ;
        RECT 12.600 165.800 13.000 166.200 ;
        RECT 9.400 164.800 9.800 165.200 ;
        RECT 12.600 161.200 12.900 165.800 ;
        RECT 13.400 163.100 13.800 168.900 ;
        RECT 15.000 168.800 16.200 169.100 ;
        RECT 16.600 165.100 17.000 167.900 ;
        RECT 18.200 163.100 18.600 168.900 ;
        RECT 20.600 165.800 21.000 166.200 ;
        RECT 22.200 165.800 22.600 166.200 ;
        RECT 15.000 161.800 15.400 162.200 ;
        RECT 6.200 160.800 6.600 161.200 ;
        RECT 12.600 160.800 13.000 161.200 ;
        RECT 6.200 155.200 6.500 160.800 ;
        RECT 3.800 154.800 4.200 155.200 ;
        RECT 5.400 154.800 5.800 155.200 ;
        RECT 6.200 154.800 6.600 155.200 ;
        RECT 3.800 154.200 4.100 154.800 ;
        RECT 3.800 153.800 4.200 154.200 ;
        RECT 0.600 145.100 1.000 147.900 ;
        RECT 2.200 143.100 2.600 148.900 ;
        RECT 6.200 146.200 6.500 154.800 ;
        RECT 7.000 152.100 7.400 157.900 ;
        RECT 10.200 156.800 10.600 157.200 ;
        RECT 10.200 153.200 10.500 156.800 ;
        RECT 15.000 155.200 15.300 161.800 ;
        RECT 20.600 159.200 20.900 165.800 ;
        RECT 22.200 161.200 22.500 165.800 ;
        RECT 23.000 163.100 23.400 168.900 ;
        RECT 28.600 163.100 29.000 168.900 ;
        RECT 31.800 168.800 32.200 169.200 ;
        RECT 25.400 161.800 25.800 162.200 ;
        RECT 26.200 161.800 26.600 162.200 ;
        RECT 22.200 160.800 22.600 161.200 ;
        RECT 20.600 158.800 21.000 159.200 ;
        RECT 18.200 156.100 18.600 156.200 ;
        RECT 19.000 156.100 19.400 156.200 ;
        RECT 18.200 155.800 19.400 156.100 ;
        RECT 15.000 154.800 15.400 155.200 ;
        RECT 15.800 154.800 16.200 155.200 ;
        RECT 19.000 154.800 19.400 155.200 ;
        RECT 19.800 155.100 20.200 155.200 ;
        RECT 20.600 155.100 21.000 155.200 ;
        RECT 19.800 154.800 21.000 155.100 ;
        RECT 22.200 154.800 22.600 155.200 ;
        RECT 11.800 154.100 12.200 154.200 ;
        RECT 12.600 154.100 13.000 154.200 ;
        RECT 11.800 153.800 13.000 154.100 ;
        RECT 10.200 153.100 10.600 153.200 ;
        RECT 11.000 153.100 11.400 153.200 ;
        RECT 10.200 152.800 11.400 153.100 ;
        RECT 3.800 146.100 4.200 146.200 ;
        RECT 4.600 146.100 5.000 146.200 ;
        RECT 3.800 145.800 5.000 146.100 ;
        RECT 6.200 145.800 6.600 146.200 ;
        RECT 0.600 133.100 1.000 135.900 ;
        RECT 2.200 132.100 2.600 137.900 ;
        RECT 6.200 135.200 6.500 145.800 ;
        RECT 7.000 143.100 7.400 148.900 ;
        RECT 9.400 148.800 9.800 149.200 ;
        RECT 9.400 148.200 9.700 148.800 ;
        RECT 9.400 147.800 9.800 148.200 ;
        RECT 10.200 148.100 10.600 148.200 ;
        RECT 11.000 148.100 11.400 148.200 ;
        RECT 10.200 147.800 11.400 148.100 ;
        RECT 11.800 146.800 12.200 147.200 ;
        RECT 12.600 146.800 13.000 147.200 ;
        RECT 13.400 147.100 13.800 147.200 ;
        RECT 14.200 147.100 14.600 147.200 ;
        RECT 13.400 146.800 14.600 147.100 ;
        RECT 11.800 146.200 12.100 146.800 ;
        RECT 12.600 146.200 12.900 146.800 ;
        RECT 15.000 146.200 15.300 154.800 ;
        RECT 15.800 154.200 16.100 154.800 ;
        RECT 19.000 154.200 19.300 154.800 ;
        RECT 15.800 153.800 16.200 154.200 ;
        RECT 16.600 153.800 17.000 154.200 ;
        RECT 19.000 153.800 19.400 154.200 ;
        RECT 16.600 153.200 16.900 153.800 ;
        RECT 16.600 152.800 17.000 153.200 ;
        RECT 18.200 151.800 18.600 152.200 ;
        RECT 15.800 147.800 16.200 148.200 ;
        RECT 15.800 147.200 16.100 147.800 ;
        RECT 15.800 146.800 16.200 147.200 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 12.600 145.800 13.000 146.200 ;
        RECT 15.000 145.800 15.400 146.200 ;
        RECT 3.000 134.700 3.400 135.100 ;
        RECT 6.200 134.800 6.600 135.200 ;
        RECT 3.000 129.200 3.300 134.700 ;
        RECT 6.200 134.200 6.500 134.800 ;
        RECT 6.200 133.800 6.600 134.200 ;
        RECT 4.600 131.800 5.000 132.200 ;
        RECT 7.000 132.100 7.400 137.900 ;
        RECT 10.200 133.100 10.600 135.900 ;
        RECT 11.000 134.800 11.400 135.200 ;
        RECT 11.000 134.200 11.300 134.800 ;
        RECT 11.000 133.800 11.400 134.200 ;
        RECT 9.400 131.800 9.800 132.200 ;
        RECT 11.800 132.100 12.200 137.900 ;
        RECT 15.000 136.200 15.300 145.800 ;
        RECT 17.400 144.800 17.800 145.200 ;
        RECT 17.400 144.200 17.700 144.800 ;
        RECT 18.200 144.200 18.500 151.800 ;
        RECT 19.800 148.100 20.200 148.200 ;
        RECT 20.600 148.100 21.000 148.200 ;
        RECT 19.800 147.800 21.000 148.100 ;
        RECT 22.200 146.200 22.500 154.800 ;
        RECT 25.400 154.200 25.700 161.800 ;
        RECT 26.200 159.200 26.500 161.800 ;
        RECT 28.600 160.800 29.000 161.200 ;
        RECT 28.600 159.200 28.900 160.800 ;
        RECT 26.200 158.800 26.600 159.200 ;
        RECT 28.600 158.800 29.000 159.200 ;
        RECT 26.200 156.100 26.600 156.200 ;
        RECT 27.000 156.100 27.400 156.200 ;
        RECT 26.200 155.800 27.400 156.100 ;
        RECT 25.400 153.800 25.800 154.200 ;
        RECT 27.000 151.800 27.400 152.200 ;
        RECT 25.400 146.800 25.800 147.200 ;
        RECT 25.400 146.200 25.700 146.800 ;
        RECT 19.000 145.800 19.400 146.200 ;
        RECT 21.400 145.800 21.800 146.200 ;
        RECT 22.200 145.800 22.600 146.200 ;
        RECT 25.400 145.800 25.800 146.200 ;
        RECT 19.000 145.200 19.300 145.800 ;
        RECT 19.000 144.800 19.400 145.200 ;
        RECT 17.400 143.800 17.800 144.200 ;
        RECT 18.200 143.800 18.600 144.200 ;
        RECT 15.000 135.800 15.400 136.200 ;
        RECT 13.400 135.100 13.800 135.200 ;
        RECT 14.200 135.100 14.600 135.200 ;
        RECT 13.400 134.800 14.600 135.100 ;
        RECT 15.800 133.800 16.200 134.200 ;
        RECT 3.000 128.800 3.400 129.200 ;
        RECT 4.600 126.200 4.900 131.800 ;
        RECT 9.400 131.200 9.700 131.800 ;
        RECT 6.200 130.800 6.600 131.200 ;
        RECT 9.400 130.800 9.800 131.200 ;
        RECT 6.200 128.200 6.500 130.800 ;
        RECT 6.200 127.800 6.600 128.200 ;
        RECT 11.800 128.100 12.200 128.200 ;
        RECT 12.600 128.100 13.000 128.200 ;
        RECT 11.800 127.800 13.000 128.100 ;
        RECT 11.000 126.800 11.400 127.200 ;
        RECT 12.600 126.800 13.000 127.200 ;
        RECT 11.000 126.200 11.300 126.800 ;
        RECT 1.400 126.100 1.800 126.200 ;
        RECT 2.200 126.100 2.600 126.200 ;
        RECT 1.400 125.800 2.600 126.100 ;
        RECT 3.800 125.800 4.200 126.200 ;
        RECT 4.600 125.800 5.000 126.200 ;
        RECT 5.400 126.100 5.800 126.200 ;
        RECT 6.200 126.100 6.600 126.200 ;
        RECT 5.400 125.800 6.600 126.100 ;
        RECT 7.000 125.800 7.400 126.200 ;
        RECT 7.800 125.800 8.200 126.200 ;
        RECT 11.000 125.800 11.400 126.200 ;
        RECT 3.800 125.200 4.100 125.800 ;
        RECT 3.800 124.800 4.200 125.200 ;
        RECT 4.600 123.800 5.000 124.200 ;
        RECT 2.200 117.100 2.600 117.200 ;
        RECT 3.000 117.100 3.400 117.200 ;
        RECT 2.200 116.800 3.400 117.100 ;
        RECT 3.800 115.800 4.200 116.200 ;
        RECT 3.800 115.200 4.100 115.800 ;
        RECT 4.600 115.200 4.900 123.800 ;
        RECT 7.000 119.200 7.300 125.800 ;
        RECT 7.000 118.800 7.400 119.200 ;
        RECT 7.800 116.200 8.100 125.800 ;
        RECT 10.200 124.800 10.600 125.200 ;
        RECT 1.400 115.100 1.800 115.200 ;
        RECT 2.200 115.100 2.600 115.200 ;
        RECT 1.400 114.800 2.600 115.100 ;
        RECT 3.800 114.800 4.200 115.200 ;
        RECT 4.600 114.800 5.000 115.200 ;
        RECT 5.400 115.100 5.800 115.200 ;
        RECT 6.200 115.100 6.600 115.200 ;
        RECT 5.400 114.800 6.600 115.100 ;
        RECT 0.600 105.100 1.000 107.900 ;
        RECT 2.200 103.100 2.600 108.900 ;
        RECT 3.800 105.800 4.200 106.200 ;
        RECT 3.800 105.200 4.100 105.800 ;
        RECT 3.800 104.800 4.200 105.200 ;
        RECT 0.600 93.100 1.000 95.900 ;
        RECT 2.200 92.100 2.600 97.900 ;
        RECT 3.000 95.100 3.400 95.200 ;
        RECT 3.800 95.100 4.200 95.200 ;
        RECT 3.000 94.800 4.200 95.100 ;
        RECT 3.000 92.800 3.400 93.200 ;
        RECT 0.600 85.100 1.000 87.900 ;
        RECT 2.200 83.100 2.600 88.900 ;
        RECT 3.000 88.200 3.300 92.800 ;
        RECT 3.000 87.800 3.400 88.200 ;
        RECT 3.000 86.100 3.400 86.200 ;
        RECT 3.800 86.100 4.200 86.200 ;
        RECT 3.000 85.800 4.200 86.100 ;
        RECT 0.600 73.100 1.000 75.900 ;
        RECT 2.200 72.100 2.600 77.900 ;
        RECT 3.000 75.100 3.400 75.200 ;
        RECT 3.800 75.100 4.200 75.200 ;
        RECT 3.000 74.800 4.200 75.100 ;
        RECT 3.800 72.800 4.200 73.200 ;
        RECT 3.000 61.800 3.400 62.200 ;
        RECT 1.400 55.100 1.800 55.200 ;
        RECT 2.200 55.100 2.600 55.200 ;
        RECT 1.400 54.800 2.600 55.100 ;
        RECT 3.000 54.200 3.300 61.800 ;
        RECT 3.800 55.200 4.100 72.800 ;
        RECT 4.600 66.200 4.900 114.800 ;
        RECT 6.200 113.800 6.600 114.200 ;
        RECT 6.200 113.200 6.500 113.800 ;
        RECT 6.200 112.800 6.600 113.200 ;
        RECT 7.000 113.100 7.400 115.900 ;
        RECT 7.800 115.800 8.200 116.200 ;
        RECT 8.600 112.100 9.000 117.900 ;
        RECT 9.400 116.800 9.800 117.200 ;
        RECT 9.400 115.100 9.700 116.800 ;
        RECT 9.400 114.700 9.800 115.100 ;
        RECT 6.200 108.800 6.600 109.200 ;
        RECT 6.200 106.200 6.500 108.800 ;
        RECT 6.200 105.800 6.600 106.200 ;
        RECT 7.000 103.100 7.400 108.900 ;
        RECT 10.200 106.200 10.500 124.800 ;
        RECT 12.600 115.200 12.900 126.800 ;
        RECT 13.400 125.100 13.800 127.900 ;
        RECT 15.000 123.100 15.400 128.900 ;
        RECT 15.800 128.200 16.100 133.800 ;
        RECT 16.600 132.100 17.000 137.900 ;
        RECT 19.000 137.100 19.400 137.200 ;
        RECT 19.800 137.100 20.200 137.200 ;
        RECT 19.000 136.800 20.200 137.100 ;
        RECT 20.600 135.800 21.000 136.200 ;
        RECT 20.600 135.200 20.900 135.800 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 20.600 134.800 21.000 135.200 ;
        RECT 19.800 132.200 20.100 134.800 ;
        RECT 19.800 131.800 20.200 132.200 ;
        RECT 15.800 127.800 16.200 128.200 ;
        RECT 15.800 125.900 16.200 126.300 ;
        RECT 15.800 125.200 16.100 125.900 ;
        RECT 15.800 124.800 16.200 125.200 ;
        RECT 19.800 123.100 20.200 128.900 ;
        RECT 21.400 125.200 21.700 145.800 ;
        RECT 22.200 136.200 22.500 145.800 ;
        RECT 27.000 138.200 27.300 151.800 ;
        RECT 28.600 144.800 29.000 145.200 ;
        RECT 27.800 141.800 28.200 142.200 ;
        RECT 27.000 137.800 27.400 138.200 ;
        RECT 25.400 136.800 25.800 137.200 ;
        RECT 26.200 136.800 26.600 137.200 ;
        RECT 25.400 136.200 25.700 136.800 ;
        RECT 22.200 135.800 22.600 136.200 ;
        RECT 25.400 135.800 25.800 136.200 ;
        RECT 22.200 135.100 22.600 135.200 ;
        RECT 23.000 135.100 23.400 135.200 ;
        RECT 22.200 134.800 23.400 135.100 ;
        RECT 23.800 134.800 24.200 135.200 ;
        RECT 23.000 130.800 23.400 131.200 ;
        RECT 22.200 128.800 22.600 129.200 ;
        RECT 22.200 128.200 22.500 128.800 ;
        RECT 22.200 127.800 22.600 128.200 ;
        RECT 23.000 125.200 23.300 130.800 ;
        RECT 23.800 126.200 24.100 134.800 ;
        RECT 25.400 133.200 25.700 135.800 ;
        RECT 25.400 132.800 25.800 133.200 ;
        RECT 26.200 132.100 26.500 136.800 ;
        RECT 27.800 136.200 28.100 141.800 ;
        RECT 28.600 139.200 28.900 144.800 ;
        RECT 30.200 143.100 30.600 148.900 ;
        RECT 28.600 138.800 29.000 139.200 ;
        RECT 31.800 136.200 32.100 168.800 ;
        RECT 32.600 165.900 33.000 166.300 ;
        RECT 32.600 158.200 32.900 165.900 ;
        RECT 33.400 163.100 33.800 168.900 ;
        RECT 43.000 168.800 43.400 169.200 ;
        RECT 51.800 169.100 52.200 169.200 ;
        RECT 52.600 169.100 53.000 169.200 ;
        RECT 43.000 168.200 43.300 168.800 ;
        RECT 34.200 167.800 34.600 168.200 ;
        RECT 34.200 167.200 34.500 167.800 ;
        RECT 34.200 166.800 34.600 167.200 ;
        RECT 35.000 165.100 35.400 167.900 ;
        RECT 43.000 167.800 43.400 168.200 ;
        RECT 41.400 166.800 41.800 167.200 ;
        RECT 42.200 166.800 42.600 167.200 ;
        RECT 41.400 166.200 41.700 166.800 ;
        RECT 36.600 166.100 37.000 166.200 ;
        RECT 37.400 166.100 37.800 166.200 ;
        RECT 36.600 165.800 37.800 166.100 ;
        RECT 38.200 165.800 38.600 166.200 ;
        RECT 41.400 165.800 41.800 166.200 ;
        RECT 38.200 164.200 38.500 165.800 ;
        RECT 38.200 163.800 38.600 164.200 ;
        RECT 32.600 157.800 33.000 158.200 ;
        RECT 35.800 153.800 36.200 154.200 ;
        RECT 32.600 146.100 33.000 146.200 ;
        RECT 33.400 146.100 33.800 146.200 ;
        RECT 32.600 145.800 33.800 146.100 ;
        RECT 35.000 143.100 35.400 148.900 ;
        RECT 35.800 147.200 36.100 153.800 ;
        RECT 36.600 153.100 37.000 155.900 ;
        RECT 38.200 152.100 38.600 157.900 ;
        RECT 42.200 155.200 42.500 166.800 ;
        RECT 43.800 165.100 44.200 167.900 ;
        RECT 45.400 163.100 45.800 168.900 ;
        RECT 49.400 166.800 49.800 167.200 ;
        RECT 46.200 165.900 46.600 166.300 ;
        RECT 49.400 166.200 49.700 166.800 ;
        RECT 46.200 165.200 46.500 165.900 ;
        RECT 49.400 165.800 49.800 166.200 ;
        RECT 46.200 164.800 46.600 165.200 ;
        RECT 50.200 163.100 50.600 168.900 ;
        RECT 51.800 168.800 53.000 169.100 ;
        RECT 53.400 166.100 53.800 166.200 ;
        RECT 54.200 166.100 54.600 166.200 ;
        RECT 53.400 165.800 54.600 166.100 ;
        RECT 60.600 165.100 61.000 167.900 ;
        RECT 61.400 166.800 61.800 167.200 ;
        RECT 61.400 166.200 61.700 166.800 ;
        RECT 61.400 165.800 61.800 166.200 ;
        RECT 62.200 163.100 62.600 168.900 ;
        RECT 63.800 165.800 64.200 166.200 ;
        RECT 63.800 159.200 64.100 165.800 ;
        RECT 67.000 163.100 67.400 168.900 ;
        RECT 80.600 165.800 81.000 166.200 ;
        RECT 87.800 166.100 88.200 166.200 ;
        RECT 88.600 166.100 89.000 166.200 ;
        RECT 87.800 165.800 89.000 166.100 ;
        RECT 80.600 165.200 80.900 165.800 ;
        RECT 80.600 164.800 81.000 165.200 ;
        RECT 87.800 164.200 88.100 165.800 ;
        RECT 91.000 165.100 91.400 167.900 ;
        RECT 91.800 166.800 92.200 167.200 ;
        RECT 91.800 165.200 92.100 166.800 ;
        RECT 91.800 164.800 92.200 165.200 ;
        RECT 67.800 163.800 68.200 164.200 ;
        RECT 87.800 163.800 88.200 164.200 ;
        RECT 57.400 158.800 57.800 159.200 ;
        RECT 63.800 158.800 64.200 159.200 ;
        RECT 53.400 158.100 53.800 158.200 ;
        RECT 54.200 158.100 54.600 158.200 ;
        RECT 39.800 154.800 40.200 155.200 ;
        RECT 42.200 154.800 42.600 155.200 ;
        RECT 39.800 152.200 40.100 154.800 ;
        RECT 39.800 151.800 40.200 152.200 ;
        RECT 42.200 150.200 42.500 154.800 ;
        RECT 43.000 152.100 43.400 157.900 ;
        RECT 53.400 157.800 54.600 158.100 ;
        RECT 47.800 154.800 48.200 155.200 ;
        RECT 51.000 154.800 51.400 155.200 ;
        RECT 51.800 154.800 52.200 155.200 ;
        RECT 52.600 154.800 53.000 155.200 ;
        RECT 47.800 154.200 48.100 154.800 ;
        RECT 47.800 153.800 48.200 154.200 ;
        RECT 49.400 154.100 49.800 154.200 ;
        RECT 50.200 154.100 50.600 154.200 ;
        RECT 49.400 153.800 50.600 154.100 ;
        RECT 45.400 152.100 45.800 152.200 ;
        RECT 44.600 151.800 45.800 152.100 ;
        RECT 42.200 149.800 42.600 150.200 ;
        RECT 43.000 149.800 43.400 150.200 ;
        RECT 35.800 146.800 36.200 147.200 ;
        RECT 36.600 145.100 37.000 147.900 ;
        RECT 39.800 147.100 40.200 147.200 ;
        RECT 40.600 147.100 41.000 147.200 ;
        RECT 39.800 146.800 41.000 147.100 ;
        RECT 42.200 146.800 42.600 147.200 ;
        RECT 42.200 146.200 42.500 146.800 ;
        RECT 39.000 145.800 39.400 146.200 ;
        RECT 42.200 145.800 42.600 146.200 ;
        RECT 39.000 143.200 39.300 145.800 ;
        RECT 41.400 145.100 41.800 145.200 ;
        RECT 42.200 145.100 42.600 145.200 ;
        RECT 41.400 144.800 42.600 145.100 ;
        RECT 39.000 142.800 39.400 143.200 ;
        RECT 42.200 142.800 42.600 143.200 ;
        RECT 40.600 138.800 41.000 139.200 ;
        RECT 36.600 137.800 37.000 138.200 ;
        RECT 36.600 137.200 36.900 137.800 ;
        RECT 33.400 137.100 33.800 137.200 ;
        RECT 34.200 137.100 34.600 137.200 ;
        RECT 33.400 136.800 34.600 137.100 ;
        RECT 36.600 136.800 37.000 137.200 ;
        RECT 27.800 135.800 28.200 136.200 ;
        RECT 29.400 135.800 29.800 136.200 ;
        RECT 30.200 136.100 30.600 136.200 ;
        RECT 31.000 136.100 31.400 136.200 ;
        RECT 30.200 135.800 31.400 136.100 ;
        RECT 31.800 135.800 32.200 136.200 ;
        RECT 27.000 135.100 27.400 135.200 ;
        RECT 27.800 135.100 28.200 135.200 ;
        RECT 27.000 134.800 28.200 135.100 ;
        RECT 29.400 134.200 29.700 135.800 ;
        RECT 31.000 134.800 31.400 135.200 ;
        RECT 32.600 135.100 33.000 135.200 ;
        RECT 33.400 135.100 33.800 135.200 ;
        RECT 32.600 134.800 33.800 135.100 ;
        RECT 35.800 134.800 36.200 135.200 ;
        RECT 31.000 134.200 31.300 134.800 ;
        RECT 35.800 134.200 36.100 134.800 ;
        RECT 29.400 133.800 29.800 134.200 ;
        RECT 31.000 133.800 31.400 134.200 ;
        RECT 35.800 133.800 36.200 134.200 ;
        RECT 38.200 133.100 38.600 133.200 ;
        RECT 39.000 133.100 39.400 133.200 ;
        RECT 39.800 133.100 40.200 135.900 ;
        RECT 38.200 132.800 39.400 133.100 ;
        RECT 25.400 131.800 26.500 132.100 ;
        RECT 37.400 131.800 37.800 132.200 ;
        RECT 23.800 125.800 24.200 126.200 ;
        RECT 20.600 124.800 21.000 125.200 ;
        RECT 21.400 124.800 21.800 125.200 ;
        RECT 23.000 124.800 23.400 125.200 ;
        RECT 12.600 114.800 13.000 115.200 ;
        RECT 12.600 109.200 12.900 114.800 ;
        RECT 13.400 112.100 13.800 117.900 ;
        RECT 15.800 116.800 16.200 117.200 ;
        RECT 15.800 115.200 16.100 116.800 ;
        RECT 16.600 115.800 17.000 116.200 ;
        RECT 16.600 115.200 16.900 115.800 ;
        RECT 15.800 114.800 16.200 115.200 ;
        RECT 16.600 114.800 17.000 115.200 ;
        RECT 19.800 114.800 20.200 115.200 ;
        RECT 15.800 113.200 16.100 114.800 ;
        RECT 19.800 114.200 20.100 114.800 ;
        RECT 17.400 114.100 17.800 114.200 ;
        RECT 18.200 114.100 18.600 114.200 ;
        RECT 17.400 113.800 18.600 114.100 ;
        RECT 19.800 113.800 20.200 114.200 ;
        RECT 15.800 112.800 16.200 113.200 ;
        RECT 18.200 111.800 18.600 112.200 ;
        RECT 12.600 108.800 13.000 109.200 ;
        RECT 16.600 108.800 17.000 109.200 ;
        RECT 15.000 107.800 15.400 108.200 ;
        RECT 11.000 107.100 11.400 107.200 ;
        RECT 11.800 107.100 12.200 107.200 ;
        RECT 11.000 106.800 12.200 107.100 ;
        RECT 13.400 106.800 13.800 107.200 ;
        RECT 13.400 106.200 13.700 106.800 ;
        RECT 10.200 105.800 10.600 106.200 ;
        RECT 11.800 106.100 12.200 106.200 ;
        RECT 12.600 106.100 13.000 106.200 ;
        RECT 11.800 105.800 13.000 106.100 ;
        RECT 13.400 105.800 13.800 106.200 ;
        RECT 9.400 102.800 9.800 103.200 ;
        RECT 9.400 102.200 9.700 102.800 ;
        RECT 9.400 101.800 9.800 102.200 ;
        RECT 7.000 92.100 7.400 97.900 ;
        RECT 9.400 97.800 9.800 98.200 ;
        RECT 9.400 97.200 9.700 97.800 ;
        RECT 9.400 96.800 9.800 97.200 ;
        RECT 10.200 94.200 10.500 105.800 ;
        RECT 13.400 98.200 13.700 105.800 ;
        RECT 15.000 102.200 15.300 107.800 ;
        RECT 15.800 105.100 16.200 107.900 ;
        RECT 16.600 107.200 16.900 108.800 ;
        RECT 16.600 106.800 17.000 107.200 ;
        RECT 17.400 103.100 17.800 108.900 ;
        RECT 18.200 106.300 18.500 111.800 ;
        RECT 19.800 107.200 20.100 113.800 ;
        RECT 20.600 108.200 20.900 124.800 ;
        RECT 25.400 124.200 25.700 131.800 ;
        RECT 35.000 129.100 35.400 129.200 ;
        RECT 35.800 129.100 36.200 129.200 ;
        RECT 26.200 125.100 26.600 127.900 ;
        RECT 27.000 126.800 27.400 127.200 ;
        RECT 24.600 124.100 25.000 124.200 ;
        RECT 25.400 124.100 25.800 124.200 ;
        RECT 24.600 123.800 25.800 124.100 ;
        RECT 25.400 121.800 25.800 122.200 ;
        RECT 25.400 118.200 25.700 121.800 ;
        RECT 21.400 112.800 21.800 113.200 ;
        RECT 22.200 113.100 22.600 115.900 ;
        RECT 21.400 108.200 21.700 112.800 ;
        RECT 23.000 111.800 23.400 112.200 ;
        RECT 23.800 112.100 24.200 117.900 ;
        RECT 25.400 117.800 25.800 118.200 ;
        RECT 27.000 115.200 27.300 126.800 ;
        RECT 27.800 123.100 28.200 128.900 ;
        RECT 29.400 126.800 29.800 127.200 ;
        RECT 29.400 126.200 29.700 126.800 ;
        RECT 29.400 125.800 29.800 126.200 ;
        RECT 32.600 123.100 33.000 128.900 ;
        RECT 35.000 128.800 36.200 129.100 ;
        RECT 35.000 127.800 35.400 128.200 ;
        RECT 25.400 114.800 25.800 115.200 ;
        RECT 27.000 114.800 27.400 115.200 ;
        RECT 25.400 113.200 25.700 114.800 ;
        RECT 24.600 112.800 25.000 113.200 ;
        RECT 25.400 112.800 25.800 113.200 ;
        RECT 20.600 107.800 21.000 108.200 ;
        RECT 21.400 107.800 21.800 108.200 ;
        RECT 19.800 106.800 20.200 107.200 ;
        RECT 18.200 105.900 18.600 106.300 ;
        RECT 22.200 103.100 22.600 108.900 ;
        RECT 15.000 101.800 15.400 102.200 ;
        RECT 13.400 97.800 13.800 98.200 ;
        RECT 15.000 96.200 15.300 101.800 ;
        RECT 15.800 98.800 16.200 99.200 ;
        RECT 15.000 95.800 15.400 96.200 ;
        RECT 15.800 95.200 16.100 98.800 ;
        RECT 18.200 97.800 18.600 98.200 ;
        RECT 19.800 97.800 20.200 98.200 ;
        RECT 16.600 95.800 17.000 96.200 ;
        RECT 16.600 95.200 16.900 95.800 ;
        RECT 11.800 94.800 12.200 95.200 ;
        RECT 12.600 94.800 13.000 95.200 ;
        RECT 14.200 95.100 14.600 95.200 ;
        RECT 15.000 95.100 15.400 95.200 ;
        RECT 14.200 94.800 15.400 95.100 ;
        RECT 15.800 94.800 16.200 95.200 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 11.800 94.200 12.100 94.800 ;
        RECT 10.200 93.800 10.600 94.200 ;
        RECT 11.800 93.800 12.200 94.200 ;
        RECT 11.800 89.800 12.200 90.200 ;
        RECT 9.400 89.100 9.800 89.200 ;
        RECT 10.200 89.100 10.600 89.200 ;
        RECT 6.200 85.800 6.600 86.200 ;
        RECT 6.200 75.200 6.500 85.800 ;
        RECT 7.000 83.100 7.400 88.900 ;
        RECT 9.400 88.800 10.600 89.100 ;
        RECT 10.200 88.100 10.600 88.200 ;
        RECT 11.000 88.100 11.400 88.200 ;
        RECT 10.200 87.800 11.400 88.100 ;
        RECT 11.800 87.200 12.100 89.800 ;
        RECT 10.200 86.800 10.600 87.200 ;
        RECT 11.800 86.800 12.200 87.200 ;
        RECT 10.200 86.200 10.500 86.800 ;
        RECT 12.600 86.200 12.900 94.800 ;
        RECT 17.400 93.800 17.800 94.200 ;
        RECT 15.000 88.800 15.400 89.200 ;
        RECT 15.000 88.200 15.300 88.800 ;
        RECT 17.400 88.200 17.700 93.800 ;
        RECT 18.200 89.200 18.500 97.800 ;
        RECT 19.800 95.200 20.100 97.800 ;
        RECT 19.800 94.800 20.200 95.200 ;
        RECT 20.600 95.100 21.000 95.200 ;
        RECT 21.400 95.100 21.800 95.200 ;
        RECT 20.600 94.800 21.800 95.100 ;
        RECT 20.600 93.800 21.000 94.200 ;
        RECT 20.600 93.200 20.900 93.800 ;
        RECT 20.600 92.800 21.000 93.200 ;
        RECT 19.000 91.800 19.400 92.200 ;
        RECT 18.200 88.800 18.600 89.200 ;
        RECT 13.400 88.100 13.800 88.200 ;
        RECT 14.200 88.100 14.600 88.200 ;
        RECT 13.400 87.800 14.600 88.100 ;
        RECT 15.000 87.800 15.400 88.200 ;
        RECT 17.400 87.800 17.800 88.200 ;
        RECT 17.400 86.800 17.800 87.200 ;
        RECT 17.400 86.200 17.700 86.800 ;
        RECT 10.200 85.800 10.600 86.200 ;
        RECT 12.600 85.800 13.000 86.200 ;
        RECT 17.400 85.800 17.800 86.200 ;
        RECT 12.600 81.100 12.900 85.800 ;
        RECT 17.400 85.100 17.800 85.200 ;
        RECT 18.200 85.100 18.600 85.200 ;
        RECT 17.400 84.800 18.600 85.100 ;
        RECT 11.800 80.800 12.900 81.100 ;
        RECT 18.200 81.800 18.600 82.200 ;
        RECT 6.200 74.800 6.600 75.200 ;
        RECT 6.200 72.200 6.500 74.800 ;
        RECT 6.200 71.800 6.600 72.200 ;
        RECT 7.000 72.100 7.400 77.900 ;
        RECT 9.400 73.800 9.800 74.200 ;
        RECT 9.400 72.200 9.700 73.800 ;
        RECT 11.800 73.200 12.100 80.800 ;
        RECT 12.600 77.800 13.000 78.200 ;
        RECT 12.600 77.200 12.900 77.800 ;
        RECT 12.600 76.800 13.000 77.200 ;
        RECT 13.400 75.800 13.800 76.200 ;
        RECT 11.000 72.800 11.400 73.200 ;
        RECT 11.800 72.800 12.200 73.200 ;
        RECT 9.400 71.800 9.800 72.200 ;
        RECT 10.200 71.800 10.600 72.200 ;
        RECT 10.200 70.200 10.500 71.800 ;
        RECT 8.600 69.800 9.000 70.200 ;
        RECT 10.200 69.800 10.600 70.200 ;
        RECT 5.400 66.800 5.800 67.200 ;
        RECT 7.800 66.800 8.200 67.200 ;
        RECT 5.400 66.200 5.700 66.800 ;
        RECT 7.800 66.200 8.100 66.800 ;
        RECT 8.600 66.200 8.900 69.800 ;
        RECT 11.000 69.200 11.300 72.800 ;
        RECT 9.400 69.100 9.800 69.200 ;
        RECT 10.200 69.100 10.600 69.200 ;
        RECT 9.400 68.800 10.600 69.100 ;
        RECT 11.000 68.800 11.400 69.200 ;
        RECT 4.600 65.800 5.000 66.200 ;
        RECT 5.400 65.800 5.800 66.200 ;
        RECT 7.800 65.800 8.200 66.200 ;
        RECT 8.600 65.800 9.000 66.200 ;
        RECT 4.600 57.200 4.900 65.800 ;
        RECT 11.800 63.100 12.200 68.900 ;
        RECT 9.400 58.800 9.800 59.200 ;
        RECT 4.600 56.800 5.000 57.200 ;
        RECT 4.600 55.200 4.900 56.800 ;
        RECT 7.000 55.800 7.400 56.200 ;
        RECT 7.000 55.200 7.300 55.800 ;
        RECT 3.800 54.800 4.200 55.200 ;
        RECT 4.600 54.800 5.000 55.200 ;
        RECT 5.400 55.100 5.800 55.200 ;
        RECT 6.200 55.100 6.600 55.200 ;
        RECT 5.400 54.800 6.600 55.100 ;
        RECT 7.000 54.800 7.400 55.200 ;
        RECT 3.000 53.800 3.400 54.200 ;
        RECT 3.000 51.800 3.400 52.200 ;
        RECT 0.600 45.100 1.000 47.900 ;
        RECT 2.200 43.100 2.600 48.900 ;
        RECT 3.000 46.300 3.300 51.800 ;
        RECT 3.000 45.900 3.400 46.300 ;
        RECT 0.600 33.100 1.000 35.900 ;
        RECT 2.200 32.100 2.600 37.900 ;
        RECT 3.800 36.200 4.100 54.800 ;
        RECT 9.400 54.200 9.700 58.800 ;
        RECT 10.200 54.800 10.600 55.200 ;
        RECT 7.800 53.800 8.200 54.200 ;
        RECT 9.400 53.800 9.800 54.200 ;
        RECT 6.200 52.800 6.600 53.200 ;
        RECT 6.200 46.200 6.500 52.800 ;
        RECT 7.800 49.200 8.100 53.800 ;
        RECT 8.600 51.800 9.000 52.200 ;
        RECT 6.200 45.800 6.600 46.200 ;
        RECT 7.000 43.100 7.400 48.900 ;
        RECT 7.800 48.800 8.200 49.200 ;
        RECT 8.600 45.200 8.900 51.800 ;
        RECT 9.400 49.800 9.800 50.200 ;
        RECT 9.400 49.200 9.700 49.800 ;
        RECT 9.400 48.800 9.800 49.200 ;
        RECT 10.200 48.200 10.500 54.800 ;
        RECT 11.000 53.100 11.400 55.900 ;
        RECT 12.600 52.100 13.000 57.900 ;
        RECT 13.400 56.200 13.700 75.800 ;
        RECT 15.800 74.800 16.200 75.200 ;
        RECT 15.800 74.200 16.100 74.800 ;
        RECT 14.200 73.800 14.600 74.200 ;
        RECT 15.800 73.800 16.200 74.200 ;
        RECT 14.200 73.200 14.500 73.800 ;
        RECT 14.200 73.100 14.600 73.200 ;
        RECT 15.000 73.100 15.400 73.200 ;
        RECT 14.200 72.800 15.400 73.100 ;
        RECT 15.800 71.800 16.200 72.200 ;
        RECT 15.800 67.200 16.100 71.800 ;
        RECT 18.200 69.200 18.500 81.800 ;
        RECT 19.000 76.200 19.300 91.800 ;
        RECT 21.400 90.200 21.700 94.800 ;
        RECT 22.200 92.800 22.600 93.200 ;
        RECT 22.200 92.200 22.500 92.800 ;
        RECT 22.200 91.800 22.600 92.200 ;
        RECT 21.400 89.800 21.800 90.200 ;
        RECT 20.600 87.800 21.000 88.200 ;
        RECT 20.600 87.200 20.900 87.800 ;
        RECT 19.800 86.800 20.200 87.200 ;
        RECT 20.600 86.800 21.000 87.200 ;
        RECT 21.400 87.100 21.800 87.200 ;
        RECT 22.200 87.100 22.600 87.200 ;
        RECT 21.400 86.800 22.600 87.100 ;
        RECT 19.800 86.200 20.100 86.800 ;
        RECT 19.800 85.800 20.200 86.200 ;
        RECT 23.000 85.200 23.300 111.800 ;
        RECT 24.600 109.200 24.900 112.800 ;
        RECT 28.600 112.100 29.000 117.900 ;
        RECT 31.800 115.800 32.200 116.200 ;
        RECT 31.800 115.200 32.100 115.800 ;
        RECT 35.000 115.200 35.300 127.800 ;
        RECT 37.400 126.200 37.700 131.800 ;
        RECT 39.000 127.800 39.400 128.200 ;
        RECT 39.000 127.200 39.300 127.800 ;
        RECT 39.000 126.800 39.400 127.200 ;
        RECT 37.400 125.800 37.800 126.200 ;
        RECT 38.200 126.100 38.600 126.200 ;
        RECT 39.000 126.100 39.400 126.200 ;
        RECT 38.200 125.800 39.400 126.100 ;
        RECT 37.400 122.200 37.700 125.800 ;
        RECT 39.800 122.800 40.200 123.200 ;
        RECT 37.400 121.800 37.800 122.200 ;
        RECT 39.800 119.200 40.100 122.800 ;
        RECT 39.800 118.800 40.200 119.200 ;
        RECT 39.800 117.800 40.200 118.200 ;
        RECT 31.800 114.800 32.200 115.200 ;
        RECT 35.000 114.800 35.400 115.200 ;
        RECT 36.600 114.800 37.000 115.200 ;
        RECT 35.000 114.200 35.300 114.800 ;
        RECT 36.600 114.200 36.900 114.800 ;
        RECT 32.600 113.800 33.000 114.200 ;
        RECT 35.000 113.800 35.400 114.200 ;
        RECT 36.600 113.800 37.000 114.200 ;
        RECT 31.000 111.800 31.400 112.200 ;
        RECT 31.000 111.200 31.300 111.800 ;
        RECT 31.000 110.800 31.400 111.200 ;
        RECT 32.600 111.100 32.900 113.800 ;
        RECT 33.400 113.100 33.800 113.200 ;
        RECT 34.200 113.100 34.600 113.200 ;
        RECT 33.400 112.800 34.600 113.100 ;
        RECT 36.600 112.800 37.000 113.200 ;
        RECT 36.600 112.200 36.900 112.800 ;
        RECT 36.600 111.800 37.000 112.200 ;
        RECT 31.800 110.800 32.900 111.100 ;
        RECT 24.600 108.800 25.000 109.200 ;
        RECT 30.200 108.800 30.600 109.200 ;
        RECT 27.800 107.800 28.200 108.200 ;
        RECT 27.800 107.200 28.100 107.800 ;
        RECT 26.200 106.800 26.600 107.200 ;
        RECT 27.800 106.800 28.200 107.200 ;
        RECT 26.200 105.100 26.500 106.800 ;
        RECT 28.600 105.800 29.000 106.200 ;
        RECT 26.200 104.800 27.300 105.100 ;
        RECT 23.800 95.800 24.200 96.200 ;
        RECT 23.800 95.200 24.100 95.800 ;
        RECT 23.800 94.800 24.200 95.200 ;
        RECT 24.600 94.800 25.000 95.200 ;
        RECT 25.400 94.800 25.800 95.200 ;
        RECT 24.600 94.200 24.900 94.800 ;
        RECT 25.400 94.200 25.700 94.800 ;
        RECT 24.600 93.800 25.000 94.200 ;
        RECT 25.400 93.800 25.800 94.200 ;
        RECT 24.600 93.200 24.900 93.800 ;
        RECT 24.600 92.800 25.000 93.200 ;
        RECT 25.400 92.100 25.800 92.200 ;
        RECT 26.200 92.100 26.600 92.200 ;
        RECT 25.400 91.800 26.600 92.100 ;
        RECT 25.400 88.800 25.800 89.200 ;
        RECT 25.400 88.200 25.700 88.800 ;
        RECT 27.000 88.200 27.300 104.800 ;
        RECT 27.800 103.800 28.200 104.200 ;
        RECT 27.800 103.200 28.100 103.800 ;
        RECT 27.800 102.800 28.200 103.200 ;
        RECT 28.600 102.100 28.900 105.800 ;
        RECT 29.400 105.100 29.800 107.900 ;
        RECT 30.200 107.200 30.500 108.800 ;
        RECT 30.200 106.800 30.600 107.200 ;
        RECT 31.000 103.100 31.400 108.900 ;
        RECT 27.800 101.800 28.900 102.100 ;
        RECT 25.400 87.800 25.800 88.200 ;
        RECT 27.000 87.800 27.400 88.200 ;
        RECT 25.400 86.100 25.800 86.200 ;
        RECT 26.200 86.100 26.600 86.200 ;
        RECT 25.400 85.800 26.600 86.100 ;
        RECT 27.800 85.200 28.100 101.800 ;
        RECT 28.600 92.100 29.000 97.900 ;
        RECT 30.200 95.800 30.600 96.200 ;
        RECT 30.200 95.200 30.500 95.800 ;
        RECT 29.400 94.800 29.800 95.200 ;
        RECT 30.200 94.800 30.600 95.200 ;
        RECT 28.600 88.800 29.000 89.200 ;
        RECT 28.600 86.200 28.900 88.800 ;
        RECT 29.400 87.200 29.700 94.800 ;
        RECT 31.000 93.800 31.400 94.200 ;
        RECT 30.200 87.800 30.600 88.200 ;
        RECT 29.400 86.800 29.800 87.200 ;
        RECT 28.600 85.800 29.000 86.200 ;
        RECT 23.000 84.800 23.400 85.200 ;
        RECT 26.200 84.800 26.600 85.200 ;
        RECT 27.000 85.100 27.400 85.200 ;
        RECT 27.800 85.100 28.200 85.200 ;
        RECT 27.000 84.800 28.200 85.100 ;
        RECT 21.400 83.800 21.800 84.200 ;
        RECT 21.400 79.200 21.700 83.800 ;
        RECT 22.200 81.800 22.600 82.200 ;
        RECT 21.400 78.800 21.800 79.200 ;
        RECT 22.200 78.200 22.500 81.800 ;
        RECT 19.800 77.800 20.200 78.200 ;
        RECT 22.200 77.800 22.600 78.200 ;
        RECT 19.000 75.800 19.400 76.200 ;
        RECT 19.800 75.200 20.100 77.800 ;
        RECT 23.000 77.200 23.300 84.800 ;
        RECT 23.800 84.100 24.200 84.200 ;
        RECT 24.600 84.100 25.000 84.200 ;
        RECT 23.800 83.800 25.000 84.100 ;
        RECT 25.400 83.800 25.800 84.200 ;
        RECT 25.400 79.200 25.700 83.800 ;
        RECT 26.200 79.200 26.500 84.800 ;
        RECT 30.200 84.200 30.500 87.800 ;
        RECT 30.200 83.800 30.600 84.200 ;
        RECT 27.800 82.800 28.200 83.200 ;
        RECT 27.800 82.200 28.100 82.800 ;
        RECT 27.800 81.800 28.200 82.200 ;
        RECT 25.400 78.800 25.800 79.200 ;
        RECT 26.200 78.800 26.600 79.200 ;
        RECT 23.000 76.800 23.400 77.200 ;
        RECT 23.800 77.100 24.200 77.200 ;
        RECT 24.600 77.100 25.000 77.200 ;
        RECT 23.800 76.800 25.000 77.100 ;
        RECT 21.400 76.100 21.800 76.200 ;
        RECT 22.200 76.100 22.600 76.200 ;
        RECT 21.400 75.800 22.600 76.100 ;
        RECT 23.000 75.800 23.400 76.200 ;
        RECT 23.000 75.200 23.300 75.800 ;
        RECT 19.000 74.800 19.400 75.200 ;
        RECT 19.800 74.800 20.200 75.200 ;
        RECT 23.000 74.800 23.400 75.200 ;
        RECT 23.800 74.800 24.200 75.200 ;
        RECT 19.000 74.100 19.300 74.800 ;
        RECT 19.000 73.800 20.100 74.100 ;
        RECT 15.800 66.800 16.200 67.200 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 15.000 66.100 15.400 66.200 ;
        RECT 14.200 65.800 15.400 66.100 ;
        RECT 13.400 55.800 13.800 56.200 ;
        RECT 15.800 55.100 16.100 66.800 ;
        RECT 16.600 63.100 17.000 68.900 ;
        RECT 18.200 68.800 18.600 69.200 ;
        RECT 18.200 65.100 18.600 67.900 ;
        RECT 19.800 67.200 20.100 73.800 ;
        RECT 20.600 73.800 21.000 74.200 ;
        RECT 20.600 73.200 20.900 73.800 ;
        RECT 20.600 72.800 21.000 73.200 ;
        RECT 23.800 69.200 24.100 74.800 ;
        RECT 26.200 73.100 26.600 75.900 ;
        RECT 27.800 72.100 28.200 77.900 ;
        RECT 29.400 75.100 29.800 75.200 ;
        RECT 30.200 75.100 30.600 75.200 ;
        RECT 29.400 74.800 30.600 75.100 ;
        RECT 31.000 75.100 31.300 93.800 ;
        RECT 31.800 93.200 32.100 110.800 ;
        RECT 38.200 109.100 38.600 109.200 ;
        RECT 39.000 109.100 39.400 109.200 ;
        RECT 32.600 105.800 33.000 106.200 ;
        RECT 32.600 105.200 32.900 105.800 ;
        RECT 32.600 104.800 33.000 105.200 ;
        RECT 35.800 103.100 36.200 108.900 ;
        RECT 38.200 108.800 39.400 109.100 ;
        RECT 39.800 106.200 40.100 117.800 ;
        RECT 40.600 116.200 40.900 138.800 ;
        RECT 41.400 132.100 41.800 137.900 ;
        RECT 41.400 121.800 41.800 122.200 ;
        RECT 40.600 115.800 41.000 116.200 ;
        RECT 39.800 105.800 40.200 106.200 ;
        RECT 32.600 101.800 33.000 102.200 ;
        RECT 31.800 92.800 32.200 93.200 ;
        RECT 31.800 86.100 32.200 86.200 ;
        RECT 32.600 86.100 32.900 101.800 ;
        RECT 33.400 92.100 33.800 97.900 ;
        RECT 35.800 96.800 36.200 97.200 ;
        RECT 37.400 97.100 37.800 97.200 ;
        RECT 38.200 97.100 38.600 97.200 ;
        RECT 37.400 96.800 38.600 97.100 ;
        RECT 35.800 96.200 36.100 96.800 ;
        RECT 35.000 93.100 35.400 95.900 ;
        RECT 35.800 95.800 36.200 96.200 ;
        RECT 36.600 95.800 37.000 96.200 ;
        RECT 36.600 95.200 36.900 95.800 ;
        RECT 36.600 94.800 37.000 95.200 ;
        RECT 36.600 91.800 37.000 92.200 ;
        RECT 31.800 85.800 32.900 86.100 ;
        RECT 33.400 86.100 33.800 86.200 ;
        RECT 33.400 85.900 34.500 86.100 ;
        RECT 33.400 85.800 34.600 85.900 ;
        RECT 34.200 85.500 34.600 85.800 ;
        RECT 35.000 85.800 35.400 86.200 ;
        RECT 35.000 85.200 35.300 85.800 ;
        RECT 35.000 84.800 35.400 85.200 ;
        RECT 36.600 84.200 36.900 91.800 ;
        RECT 37.400 90.800 37.800 91.200 ;
        RECT 37.400 86.200 37.700 90.800 ;
        RECT 39.000 86.800 39.400 87.200 ;
        RECT 37.400 85.800 37.800 86.200 ;
        RECT 39.000 84.200 39.300 86.800 ;
        RECT 35.000 83.800 35.400 84.200 ;
        RECT 36.600 83.800 37.000 84.200 ;
        RECT 39.000 83.800 39.400 84.200 ;
        RECT 35.000 79.200 35.300 83.800 ;
        RECT 39.800 82.200 40.100 105.800 ;
        RECT 40.600 104.200 40.900 115.800 ;
        RECT 41.400 115.200 41.700 121.800 ;
        RECT 42.200 115.200 42.500 142.800 ;
        RECT 43.000 134.200 43.300 149.800 ;
        RECT 43.800 148.800 44.200 149.200 ;
        RECT 43.800 148.200 44.100 148.800 ;
        RECT 43.800 147.800 44.200 148.200 ;
        RECT 44.600 147.200 44.900 151.800 ;
        RECT 44.600 146.800 45.000 147.200 ;
        RECT 46.200 144.800 46.600 145.200 ;
        RECT 47.000 145.100 47.400 147.900 ;
        RECT 47.800 147.200 48.100 153.800 ;
        RECT 49.400 152.100 49.800 152.200 ;
        RECT 50.200 152.100 50.600 152.200 ;
        RECT 49.400 151.800 50.600 152.100 ;
        RECT 51.000 151.200 51.300 154.800 ;
        RECT 51.800 153.200 52.100 154.800 ;
        RECT 51.800 152.800 52.200 153.200 ;
        RECT 51.000 150.800 51.400 151.200 ;
        RECT 51.800 150.200 52.100 152.800 ;
        RECT 49.400 149.800 49.800 150.200 ;
        RECT 51.800 149.800 52.200 150.200 ;
        RECT 47.800 146.800 48.200 147.200 ;
        RECT 46.200 144.200 46.500 144.800 ;
        RECT 46.200 143.800 46.600 144.200 ;
        RECT 45.400 141.800 45.800 142.200 ;
        RECT 43.800 134.800 44.200 135.200 ;
        RECT 43.000 133.800 43.400 134.200 ;
        RECT 43.000 133.200 43.300 133.800 ;
        RECT 43.000 132.800 43.400 133.200 ;
        RECT 43.000 128.800 43.400 129.200 ;
        RECT 43.000 128.200 43.300 128.800 ;
        RECT 43.000 127.800 43.400 128.200 ;
        RECT 43.800 127.200 44.100 134.800 ;
        RECT 45.400 131.200 45.700 141.800 ;
        RECT 46.200 132.100 46.600 137.900 ;
        RECT 47.800 135.200 48.100 146.800 ;
        RECT 48.600 143.100 49.000 148.900 ;
        RECT 49.400 148.200 49.700 149.800 ;
        RECT 49.400 147.800 49.800 148.200 ;
        RECT 49.400 146.800 49.800 147.200 ;
        RECT 49.400 146.300 49.700 146.800 ;
        RECT 49.400 145.900 49.800 146.300 ;
        RECT 52.600 146.200 52.900 154.800 ;
        RECT 57.400 154.200 57.700 158.800 ;
        RECT 59.800 156.100 60.200 156.200 ;
        RECT 60.600 156.100 61.000 156.200 ;
        RECT 59.800 155.800 61.000 156.100 ;
        RECT 67.800 155.200 68.100 163.800 ;
        RECT 92.600 163.100 93.000 168.900 ;
        RECT 94.200 165.800 94.600 166.200 ;
        RECT 94.200 165.200 94.500 165.800 ;
        RECT 94.200 164.800 94.600 165.200 ;
        RECT 97.400 163.100 97.800 168.900 ;
        RECT 104.600 166.800 105.000 167.200 ;
        RECT 104.600 166.200 104.900 166.800 ;
        RECT 100.600 165.800 101.000 166.200 ;
        RECT 101.400 166.100 101.800 166.200 ;
        RECT 102.200 166.100 102.600 166.200 ;
        RECT 101.400 165.800 102.600 166.100 ;
        RECT 104.600 165.800 105.000 166.200 ;
        RECT 100.600 164.200 100.900 165.800 ;
        RECT 100.600 163.800 101.000 164.200 ;
        RECT 109.400 163.100 109.800 168.900 ;
        RECT 112.600 166.800 113.000 167.200 ;
        RECT 111.000 166.100 111.400 166.200 ;
        RECT 111.800 166.100 112.200 166.200 ;
        RECT 111.000 165.800 112.200 166.100 ;
        RECT 69.400 161.800 69.800 162.200 ;
        RECT 72.600 161.800 73.000 162.200 ;
        RECT 83.800 161.800 84.200 162.200 ;
        RECT 99.800 162.100 100.200 162.200 ;
        RECT 99.800 161.800 100.900 162.100 ;
        RECT 69.400 161.200 69.700 161.800 ;
        RECT 69.400 160.800 69.800 161.200 ;
        RECT 72.600 158.200 72.900 161.800 ;
        RECT 59.800 155.100 60.200 155.200 ;
        RECT 60.600 155.100 61.000 155.200 ;
        RECT 59.800 154.800 61.000 155.100 ;
        RECT 61.400 154.800 61.800 155.200 ;
        RECT 67.800 154.800 68.200 155.200 ;
        RECT 57.400 153.800 57.800 154.200 ;
        RECT 59.000 151.800 59.400 152.200 ;
        RECT 55.800 149.100 56.200 149.200 ;
        RECT 56.600 149.100 57.000 149.200 ;
        RECT 52.600 145.800 53.000 146.200 ;
        RECT 53.400 143.100 53.800 148.900 ;
        RECT 55.800 148.800 57.000 149.100 ;
        RECT 54.200 145.800 54.600 146.200 ;
        RECT 57.400 145.800 57.800 146.200 ;
        RECT 54.200 135.200 54.500 145.800 ;
        RECT 57.400 139.200 57.700 145.800 ;
        RECT 59.000 144.200 59.300 151.800 ;
        RECT 61.400 151.200 61.700 154.800 ;
        RECT 63.800 154.100 64.200 154.200 ;
        RECT 64.600 154.100 65.000 154.200 ;
        RECT 63.800 153.800 65.000 154.100 ;
        RECT 68.600 152.800 69.000 153.200 ;
        RECT 61.400 150.800 61.800 151.200 ;
        RECT 59.800 148.800 60.200 149.200 ;
        RECT 67.800 148.800 68.200 149.200 ;
        RECT 59.800 147.200 60.100 148.800 ;
        RECT 62.200 148.100 62.600 148.200 ;
        RECT 63.000 148.100 63.400 148.200 ;
        RECT 62.200 147.800 63.400 148.100 ;
        RECT 64.600 147.800 65.000 148.200 ;
        RECT 59.800 146.800 60.200 147.200 ;
        RECT 63.000 147.100 63.400 147.200 ;
        RECT 63.800 147.100 64.200 147.200 ;
        RECT 63.000 146.800 64.200 147.100 ;
        RECT 64.600 146.200 64.900 147.800 ;
        RECT 66.200 147.100 66.600 147.200 ;
        RECT 67.000 147.100 67.400 147.200 ;
        RECT 66.200 146.800 67.400 147.100 ;
        RECT 64.600 145.800 65.000 146.200 ;
        RECT 60.600 145.100 61.000 145.200 ;
        RECT 61.400 145.100 61.800 145.200 ;
        RECT 60.600 144.800 61.800 145.100 ;
        RECT 65.400 144.800 65.800 145.200 ;
        RECT 59.000 143.800 59.400 144.200 ;
        RECT 58.200 141.800 58.600 142.200 ;
        RECT 60.600 141.800 61.000 142.200 ;
        RECT 57.400 138.800 57.800 139.200 ;
        RECT 55.800 137.100 56.200 137.200 ;
        RECT 56.600 137.100 57.000 137.200 ;
        RECT 55.800 136.800 57.000 137.100 ;
        RECT 58.200 136.200 58.500 141.800 ;
        RECT 60.600 136.200 60.900 141.800 ;
        RECT 65.400 138.200 65.700 144.800 ;
        RECT 65.400 137.800 65.800 138.200 ;
        RECT 61.400 137.100 61.800 137.200 ;
        RECT 62.200 137.100 62.600 137.200 ;
        RECT 61.400 136.800 62.600 137.100 ;
        RECT 65.400 136.200 65.700 137.800 ;
        RECT 66.200 136.800 66.600 137.200 ;
        RECT 66.200 136.200 66.500 136.800 ;
        RECT 55.000 135.800 55.400 136.200 ;
        RECT 58.200 135.800 58.600 136.200 ;
        RECT 59.000 136.100 59.400 136.200 ;
        RECT 59.800 136.100 60.200 136.200 ;
        RECT 59.000 135.800 60.200 136.100 ;
        RECT 60.600 135.800 61.000 136.200 ;
        RECT 65.400 135.800 65.800 136.200 ;
        RECT 66.200 135.800 66.600 136.200 ;
        RECT 47.800 134.800 48.200 135.200 ;
        RECT 49.400 135.100 49.800 135.200 ;
        RECT 50.200 135.100 50.600 135.200 ;
        RECT 49.400 134.800 50.600 135.100 ;
        RECT 53.400 134.800 53.800 135.200 ;
        RECT 54.200 134.800 54.600 135.200 ;
        RECT 53.400 134.200 53.700 134.800 ;
        RECT 51.800 134.100 52.200 134.200 ;
        RECT 52.600 134.100 53.000 134.200 ;
        RECT 51.800 133.800 53.000 134.100 ;
        RECT 53.400 133.800 53.800 134.200 ;
        RECT 51.000 132.800 51.400 133.200 ;
        RECT 52.600 132.800 53.000 133.200 ;
        RECT 48.600 132.100 49.000 132.200 ;
        RECT 49.400 132.100 49.800 132.200 ;
        RECT 48.600 131.800 49.800 132.100 ;
        RECT 44.600 130.800 45.000 131.200 ;
        RECT 45.400 130.800 45.800 131.200 ;
        RECT 43.800 126.800 44.200 127.200 ;
        RECT 44.600 126.200 44.900 130.800 ;
        RECT 49.400 128.200 49.700 131.800 ;
        RECT 51.000 130.200 51.300 132.800 ;
        RECT 51.000 129.800 51.400 130.200 ;
        RECT 45.400 127.800 45.800 128.200 ;
        RECT 49.400 127.800 49.800 128.200 ;
        RECT 45.400 127.200 45.700 127.800 ;
        RECT 45.400 126.800 45.800 127.200 ;
        RECT 43.800 125.800 44.200 126.200 ;
        RECT 44.600 125.800 45.000 126.200 ;
        RECT 43.800 125.200 44.100 125.800 ;
        RECT 43.800 124.800 44.200 125.200 ;
        RECT 43.000 117.100 43.400 117.200 ;
        RECT 43.800 117.100 44.200 117.200 ;
        RECT 43.000 116.800 44.200 117.100 ;
        RECT 44.600 116.200 44.900 125.800 ;
        RECT 50.200 125.100 50.600 127.900 ;
        RECT 51.000 126.800 51.400 127.200 ;
        RECT 44.600 115.800 45.000 116.200 ;
        RECT 41.400 114.800 41.800 115.200 ;
        RECT 42.200 114.800 42.600 115.200 ;
        RECT 47.000 114.800 47.400 115.200 ;
        RECT 41.400 107.200 41.700 114.800 ;
        RECT 42.200 114.200 42.500 114.800 ;
        RECT 42.200 113.800 42.600 114.200 ;
        RECT 42.200 113.200 42.500 113.800 ;
        RECT 47.000 113.200 47.300 114.800 ;
        RECT 42.200 112.800 42.600 113.200 ;
        RECT 47.000 112.800 47.400 113.200 ;
        RECT 47.800 113.100 48.200 115.900 ;
        RECT 47.000 111.800 47.400 112.200 ;
        RECT 49.400 112.100 49.800 117.900 ;
        RECT 50.200 116.800 50.600 117.200 ;
        RECT 50.200 115.100 50.500 116.800 ;
        RECT 50.200 114.700 50.600 115.100 ;
        RECT 51.000 114.200 51.300 126.800 ;
        RECT 51.800 123.100 52.200 128.900 ;
        RECT 52.600 128.200 52.900 132.800 ;
        RECT 53.400 128.200 53.700 133.800 ;
        RECT 52.600 127.800 53.000 128.200 ;
        RECT 53.400 127.800 53.800 128.200 ;
        RECT 53.400 126.800 53.800 127.200 ;
        RECT 53.400 126.200 53.700 126.800 ;
        RECT 54.200 126.200 54.500 134.800 ;
        RECT 53.400 125.800 53.800 126.200 ;
        RECT 54.200 125.800 54.600 126.200 ;
        RECT 51.800 121.800 52.200 122.200 ;
        RECT 51.000 113.800 51.400 114.200 ;
        RECT 51.800 113.100 52.100 121.800 ;
        RECT 51.000 112.800 52.100 113.100 ;
        RECT 46.200 108.800 46.600 109.200 ;
        RECT 46.200 108.200 46.500 108.800 ;
        RECT 46.200 107.800 46.600 108.200 ;
        RECT 46.200 107.200 46.500 107.800 ;
        RECT 47.000 107.200 47.300 111.800 ;
        RECT 51.000 109.200 51.300 112.800 ;
        RECT 54.200 112.100 54.600 117.900 ;
        RECT 55.000 116.200 55.300 135.800 ;
        RECT 55.800 134.800 56.200 135.200 ;
        RECT 61.400 134.800 61.800 135.200 ;
        RECT 55.800 134.200 56.100 134.800 ;
        RECT 55.800 133.800 56.200 134.200 ;
        RECT 58.200 133.800 58.600 134.200 ;
        RECT 58.200 132.200 58.500 133.800 ;
        RECT 61.400 133.200 61.700 134.800 ;
        RECT 67.800 134.200 68.100 148.800 ;
        RECT 68.600 143.200 68.900 152.800 ;
        RECT 69.400 152.100 69.800 157.900 ;
        RECT 72.600 157.800 73.000 158.200 ;
        RECT 70.200 155.800 70.600 156.200 ;
        RECT 70.200 155.200 70.500 155.800 ;
        RECT 70.200 154.800 70.600 155.200 ;
        RECT 72.600 154.800 73.000 155.200 ;
        RECT 72.600 154.200 72.900 154.800 ;
        RECT 72.600 153.800 73.000 154.200 ;
        RECT 73.400 152.800 73.800 153.200 ;
        RECT 73.400 151.200 73.700 152.800 ;
        RECT 74.200 152.100 74.600 157.900 ;
        RECT 75.000 153.800 75.400 154.200 ;
        RECT 73.400 150.800 73.800 151.200 ;
        RECT 68.600 142.800 69.000 143.200 ;
        RECT 71.000 143.100 71.400 148.900 ;
        RECT 68.600 140.800 69.000 141.200 ;
        RECT 68.600 134.200 68.900 140.800 ;
        RECT 70.200 138.800 70.600 139.200 ;
        RECT 70.200 136.200 70.500 138.800 ;
        RECT 70.200 135.800 70.600 136.200 ;
        RECT 71.800 135.800 72.200 136.200 ;
        RECT 71.800 135.200 72.100 135.800 ;
        RECT 73.400 135.200 73.700 150.800 ;
        RECT 75.000 148.200 75.300 153.800 ;
        RECT 75.800 153.100 76.200 155.900 ;
        RECT 76.600 154.800 77.000 155.200 ;
        RECT 79.000 154.800 79.400 155.200 ;
        RECT 76.600 154.200 76.900 154.800 ;
        RECT 79.000 154.200 79.300 154.800 ;
        RECT 76.600 153.800 77.000 154.200 ;
        RECT 77.400 154.100 77.800 154.200 ;
        RECT 77.400 153.800 78.500 154.100 ;
        RECT 79.000 153.800 79.400 154.200 ;
        RECT 75.000 147.800 75.400 148.200 ;
        RECT 75.000 145.900 75.400 146.300 ;
        RECT 75.000 139.200 75.300 145.900 ;
        RECT 75.800 143.100 76.200 148.900 ;
        RECT 77.400 145.100 77.800 147.900 ;
        RECT 78.200 146.200 78.500 153.800 ;
        RECT 79.000 152.800 79.400 153.200 ;
        RECT 79.800 153.100 80.200 155.900 ;
        RECT 80.600 155.800 81.000 156.200 ;
        RECT 80.600 154.200 80.900 155.800 ;
        RECT 80.600 153.800 81.000 154.200 ;
        RECT 79.000 149.200 79.300 152.800 ;
        RECT 81.400 152.100 81.800 157.900 ;
        RECT 82.200 155.000 82.600 155.100 ;
        RECT 83.000 155.000 83.400 155.100 ;
        RECT 82.200 154.700 83.400 155.000 ;
        RECT 80.600 149.800 81.000 150.200 ;
        RECT 79.000 148.800 79.400 149.200 ;
        RECT 79.800 147.800 80.200 148.200 ;
        RECT 78.200 145.800 78.600 146.200 ;
        RECT 75.000 138.800 75.400 139.200 ;
        RECT 77.400 138.800 77.800 139.200 ;
        RECT 77.400 136.200 77.700 138.800 ;
        RECT 75.800 135.800 76.200 136.200 ;
        RECT 77.400 135.800 77.800 136.200 ;
        RECT 75.800 135.200 76.100 135.800 ;
        RECT 78.200 135.200 78.500 145.800 ;
        RECT 79.800 145.200 80.100 147.800 ;
        RECT 80.600 146.200 80.900 149.800 ;
        RECT 83.800 146.200 84.100 161.800 ;
        RECT 92.600 159.100 93.000 159.200 ;
        RECT 93.400 159.100 93.800 159.200 ;
        RECT 92.600 158.800 93.800 159.100 ;
        RECT 86.200 152.100 86.600 157.900 ;
        RECT 90.200 155.100 90.600 155.200 ;
        RECT 91.000 155.100 91.400 155.200 ;
        RECT 90.200 154.800 91.400 155.100 ;
        RECT 91.800 154.800 92.200 155.200 ;
        RECT 91.800 153.200 92.100 154.800 ;
        RECT 100.600 153.200 100.900 161.800 ;
        RECT 107.000 161.800 107.400 162.200 ;
        RECT 101.400 156.800 101.800 157.200 ;
        RECT 105.400 156.800 105.800 157.200 ;
        RECT 101.400 156.200 101.700 156.800 ;
        RECT 101.400 155.800 101.800 156.200 ;
        RECT 101.400 155.100 101.800 155.200 ;
        RECT 102.200 155.100 102.600 155.200 ;
        RECT 101.400 154.800 102.600 155.100 ;
        RECT 103.000 154.800 103.400 155.200 ;
        RECT 91.800 152.800 92.200 153.200 ;
        RECT 96.600 152.800 97.000 153.200 ;
        RECT 97.400 152.800 97.800 153.200 ;
        RECT 100.600 152.800 101.000 153.200 ;
        RECT 96.600 152.200 96.900 152.800 ;
        RECT 97.400 152.200 97.700 152.800 ;
        RECT 88.600 152.100 89.000 152.200 ;
        RECT 87.800 151.800 89.000 152.100 ;
        RECT 96.600 151.800 97.000 152.200 ;
        RECT 97.400 151.800 97.800 152.200 ;
        RECT 84.600 146.800 85.000 147.200 ;
        RECT 84.600 146.200 84.900 146.800 ;
        RECT 80.600 145.800 81.000 146.200 ;
        RECT 81.400 146.100 81.800 146.200 ;
        RECT 82.200 146.100 82.600 146.200 ;
        RECT 81.400 145.800 82.600 146.100 ;
        RECT 83.800 145.800 84.200 146.200 ;
        RECT 84.600 145.800 85.000 146.200 ;
        RECT 87.800 145.200 88.100 151.800 ;
        RECT 98.200 149.800 98.600 150.200 ;
        RECT 79.800 144.800 80.200 145.200 ;
        RECT 81.400 144.800 81.800 145.200 ;
        RECT 87.800 144.800 88.200 145.200 ;
        RECT 80.600 142.800 81.000 143.200 ;
        RECT 79.000 141.800 79.400 142.200 ;
        RECT 71.800 134.800 72.200 135.200 ;
        RECT 72.600 134.800 73.000 135.200 ;
        RECT 73.400 134.800 73.800 135.200 ;
        RECT 75.800 134.800 76.200 135.200 ;
        RECT 78.200 134.800 78.600 135.200 ;
        RECT 72.600 134.200 72.900 134.800 ;
        RECT 63.800 133.800 64.200 134.200 ;
        RECT 67.800 133.800 68.200 134.200 ;
        RECT 68.600 133.800 69.000 134.200 ;
        RECT 72.600 133.800 73.000 134.200 ;
        RECT 61.400 132.800 61.800 133.200 ;
        RECT 58.200 131.800 58.600 132.200 ;
        RECT 59.800 131.800 60.200 132.200 ;
        RECT 59.000 129.800 59.400 130.200 ;
        RECT 59.000 129.200 59.300 129.800 ;
        RECT 56.600 123.100 57.000 128.900 ;
        RECT 59.000 128.800 59.400 129.200 ;
        RECT 59.800 126.200 60.100 131.800 ;
        RECT 60.600 127.800 61.000 128.200 ;
        RECT 60.600 127.200 60.900 127.800 ;
        RECT 61.400 127.200 61.700 132.800 ;
        RECT 62.200 131.800 62.600 132.200 ;
        RECT 60.600 126.800 61.000 127.200 ;
        RECT 61.400 126.800 61.800 127.200 ;
        RECT 59.800 125.800 60.200 126.200 ;
        RECT 60.600 126.100 61.000 126.200 ;
        RECT 61.400 126.100 61.800 126.200 ;
        RECT 60.600 125.800 61.800 126.100 ;
        RECT 62.200 125.200 62.500 131.800 ;
        RECT 63.800 130.200 64.100 133.800 ;
        RECT 67.800 133.200 68.100 133.800 ;
        RECT 67.800 132.800 68.200 133.200 ;
        RECT 71.000 133.100 71.400 133.200 ;
        RECT 71.800 133.100 72.200 133.200 ;
        RECT 71.000 132.800 72.200 133.100 ;
        RECT 73.400 132.200 73.700 134.800 ;
        RECT 79.000 134.200 79.300 141.800 ;
        RECT 79.800 137.800 80.200 138.200 ;
        RECT 79.800 136.200 80.100 137.800 ;
        RECT 79.800 135.800 80.200 136.200 ;
        RECT 80.600 135.100 80.900 142.800 ;
        RECT 79.800 134.800 80.900 135.100 ;
        RECT 79.000 133.800 79.400 134.200 ;
        RECT 64.600 131.800 65.000 132.200 ;
        RECT 67.000 131.800 67.400 132.200 ;
        RECT 70.200 131.800 70.600 132.200 ;
        RECT 73.400 131.800 73.800 132.200 ;
        RECT 77.400 131.800 77.800 132.200 ;
        RECT 63.800 129.800 64.200 130.200 ;
        RECT 63.000 128.800 63.400 129.200 ;
        RECT 63.000 125.200 63.300 128.800 ;
        RECT 63.800 126.800 64.200 127.200 ;
        RECT 63.800 126.200 64.100 126.800 ;
        RECT 63.800 125.800 64.200 126.200 ;
        RECT 64.600 125.200 64.900 131.800 ;
        RECT 67.000 130.200 67.300 131.800 ;
        RECT 70.200 131.100 70.500 131.800 ;
        RECT 70.200 130.800 71.300 131.100 ;
        RECT 67.000 129.800 67.400 130.200 ;
        RECT 70.200 129.800 70.600 130.200 ;
        RECT 67.800 126.800 68.200 127.200 ;
        RECT 68.600 126.800 69.000 127.200 ;
        RECT 67.800 126.200 68.100 126.800 ;
        RECT 65.400 126.100 65.800 126.200 ;
        RECT 66.200 126.100 66.600 126.200 ;
        RECT 65.400 125.800 66.600 126.100 ;
        RECT 67.800 125.800 68.200 126.200 ;
        RECT 68.600 125.200 68.900 126.800 ;
        RECT 70.200 126.200 70.500 129.800 ;
        RECT 70.200 125.800 70.600 126.200 ;
        RECT 62.200 124.800 62.600 125.200 ;
        RECT 63.000 124.800 63.400 125.200 ;
        RECT 64.600 124.800 65.000 125.200 ;
        RECT 68.600 124.800 69.000 125.200 ;
        RECT 71.000 124.200 71.300 130.800 ;
        RECT 75.800 128.800 76.200 129.200 ;
        RECT 75.800 128.200 76.100 128.800 ;
        RECT 75.800 127.800 76.200 128.200 ;
        RECT 76.600 126.800 77.000 127.200 ;
        RECT 72.600 126.100 73.000 126.200 ;
        RECT 73.400 126.100 73.800 126.200 ;
        RECT 72.600 125.800 73.800 126.100 ;
        RECT 71.800 125.100 72.200 125.200 ;
        RECT 72.600 125.100 73.000 125.200 ;
        RECT 71.800 124.800 73.000 125.100 ;
        RECT 74.200 124.800 74.600 125.200 ;
        RECT 74.200 124.200 74.500 124.800 ;
        RECT 60.600 123.800 61.000 124.200 ;
        RECT 63.800 124.100 64.200 124.200 ;
        RECT 64.600 124.100 65.000 124.200 ;
        RECT 63.800 123.800 65.000 124.100 ;
        RECT 66.200 124.100 66.600 124.200 ;
        RECT 67.000 124.100 67.400 124.200 ;
        RECT 66.200 123.800 67.400 124.100 ;
        RECT 71.000 123.800 71.400 124.200 ;
        RECT 74.200 123.800 74.600 124.200 ;
        RECT 60.600 123.200 60.900 123.800 ;
        RECT 60.600 122.800 61.000 123.200 ;
        RECT 72.600 122.800 73.000 123.200 ;
        RECT 71.800 121.800 72.200 122.200 ;
        RECT 56.600 116.800 57.000 117.200 ;
        RECT 55.000 115.800 55.400 116.200 ;
        RECT 56.600 115.200 56.900 116.800 ;
        RECT 56.600 114.800 57.000 115.200 ;
        RECT 57.400 111.800 57.800 112.200 ;
        RECT 59.800 112.100 60.200 117.900 ;
        RECT 63.000 114.800 63.400 115.200 ;
        RECT 54.200 109.800 54.600 110.200 ;
        RECT 54.200 109.200 54.500 109.800 ;
        RECT 51.000 108.800 51.400 109.200 ;
        RECT 54.200 108.800 54.600 109.200 ;
        RECT 57.400 108.200 57.700 111.800 ;
        RECT 63.000 111.200 63.300 114.800 ;
        RECT 64.600 112.100 65.000 117.900 ;
        RECT 71.800 117.200 72.100 121.800 ;
        RECT 71.800 116.800 72.200 117.200 ;
        RECT 65.400 113.800 65.800 114.200 ;
        RECT 65.400 113.200 65.700 113.800 ;
        RECT 65.400 112.800 65.800 113.200 ;
        RECT 66.200 113.100 66.600 115.900 ;
        RECT 72.600 115.200 72.900 122.800 ;
        RECT 76.600 122.200 76.900 126.800 ;
        RECT 77.400 125.200 77.700 131.800 ;
        RECT 79.800 129.200 80.100 134.800 ;
        RECT 81.400 134.200 81.700 144.800 ;
        RECT 91.000 143.100 91.400 148.900 ;
        RECT 92.600 147.100 93.000 147.200 ;
        RECT 93.400 147.100 93.800 147.200 ;
        RECT 92.600 146.800 93.800 147.100 ;
        RECT 93.400 146.100 93.800 146.200 ;
        RECT 94.200 146.100 94.600 146.200 ;
        RECT 93.400 145.800 94.600 146.100 ;
        RECT 95.800 143.100 96.200 148.900 ;
        RECT 97.400 145.100 97.800 147.900 ;
        RECT 98.200 145.200 98.500 149.800 ;
        RECT 99.000 148.800 99.400 149.200 ;
        RECT 99.000 148.200 99.300 148.800 ;
        RECT 99.000 147.800 99.400 148.200 ;
        RECT 99.800 146.800 100.200 147.200 ;
        RECT 99.800 146.200 100.100 146.800 ;
        RECT 100.600 146.200 100.900 152.800 ;
        RECT 102.200 150.200 102.500 154.800 ;
        RECT 103.000 154.200 103.300 154.800 ;
        RECT 103.000 153.800 103.400 154.200 ;
        RECT 103.800 151.800 104.200 152.200 ;
        RECT 104.600 151.800 105.000 152.200 ;
        RECT 101.400 149.800 101.800 150.200 ;
        RECT 102.200 149.800 102.600 150.200 ;
        RECT 101.400 149.200 101.700 149.800 ;
        RECT 101.400 148.800 101.800 149.200 ;
        RECT 101.400 147.800 101.800 148.200 ;
        RECT 101.400 147.200 101.700 147.800 ;
        RECT 101.400 146.800 101.800 147.200 ;
        RECT 99.800 145.800 100.200 146.200 ;
        RECT 100.600 145.800 101.000 146.200 ;
        RECT 98.200 144.800 98.600 145.200 ;
        RECT 87.800 142.100 88.200 142.200 ;
        RECT 88.600 142.100 89.000 142.200 ;
        RECT 87.800 141.800 89.000 142.100 ;
        RECT 93.400 141.800 93.800 142.200 ;
        RECT 91.800 136.100 92.200 136.200 ;
        RECT 92.600 136.100 93.000 136.200 ;
        RECT 91.800 135.800 93.000 136.100 ;
        RECT 84.600 135.100 85.000 135.200 ;
        RECT 85.400 135.100 85.800 135.200 ;
        RECT 84.600 134.800 85.800 135.100 ;
        RECT 87.000 135.100 87.400 135.200 ;
        RECT 87.800 135.100 88.200 135.200 ;
        RECT 87.000 134.800 88.200 135.100 ;
        RECT 92.600 134.800 93.000 135.200 ;
        RECT 81.400 133.800 81.800 134.200 ;
        RECT 83.800 133.800 84.200 134.200 ;
        RECT 87.800 133.800 88.200 134.200 ;
        RECT 82.200 133.100 82.600 133.200 ;
        RECT 83.000 133.100 83.400 133.200 ;
        RECT 82.200 132.800 83.400 133.100 ;
        RECT 80.600 131.800 81.000 132.200 ;
        RECT 79.800 128.800 80.200 129.200 ;
        RECT 78.200 126.100 78.600 126.200 ;
        RECT 79.000 126.100 79.400 126.200 ;
        RECT 78.200 125.800 79.400 126.100 ;
        RECT 77.400 124.800 77.800 125.200 ;
        RECT 75.000 121.800 75.400 122.200 ;
        RECT 76.600 121.800 77.000 122.200 ;
        RECT 74.200 116.800 74.600 117.200 ;
        RECT 71.000 115.100 71.400 115.200 ;
        RECT 71.800 115.100 72.200 115.200 ;
        RECT 71.000 114.800 72.200 115.100 ;
        RECT 72.600 114.800 73.000 115.200 ;
        RECT 67.000 112.800 67.400 113.200 ;
        RECT 69.400 112.800 69.800 113.200 ;
        RECT 59.800 110.800 60.200 111.200 ;
        RECT 63.000 110.800 63.400 111.200 ;
        RECT 59.800 109.200 60.100 110.800 ;
        RECT 59.800 108.800 60.200 109.200 ;
        RECT 67.000 109.100 67.300 112.800 ;
        RECT 67.800 109.100 68.200 109.200 ;
        RECT 67.000 108.800 68.200 109.100 ;
        RECT 55.000 107.800 55.400 108.200 ;
        RECT 55.800 107.800 56.200 108.200 ;
        RECT 57.400 108.100 57.800 108.200 ;
        RECT 58.200 108.100 58.600 108.200 ;
        RECT 57.400 107.800 58.600 108.100 ;
        RECT 55.000 107.200 55.300 107.800 ;
        RECT 41.400 106.800 41.800 107.200 ;
        RECT 46.200 106.800 46.600 107.200 ;
        RECT 47.000 106.800 47.400 107.200 ;
        RECT 52.600 107.100 53.000 107.200 ;
        RECT 53.400 107.100 53.800 107.200 ;
        RECT 52.600 106.800 53.800 107.100 ;
        RECT 55.000 106.800 55.400 107.200 ;
        RECT 55.800 106.200 56.100 107.800 ;
        RECT 67.000 107.200 67.300 108.800 ;
        RECT 57.400 106.800 57.800 107.200 ;
        RECT 60.600 106.800 61.000 107.200 ;
        RECT 65.400 106.800 65.800 107.200 ;
        RECT 67.000 106.800 67.400 107.200 ;
        RECT 41.400 106.100 41.800 106.200 ;
        RECT 42.200 106.100 42.600 106.200 ;
        RECT 50.200 106.100 50.600 106.200 ;
        RECT 41.400 105.800 42.600 106.100 ;
        RECT 49.400 105.800 50.600 106.100 ;
        RECT 52.600 105.800 53.000 106.200 ;
        RECT 55.800 105.800 56.200 106.200 ;
        RECT 56.600 105.800 57.000 106.200 ;
        RECT 43.000 104.800 43.400 105.200 ;
        RECT 47.000 105.100 47.400 105.200 ;
        RECT 47.800 105.100 48.200 105.200 ;
        RECT 47.000 104.800 48.200 105.100 ;
        RECT 48.600 104.800 49.000 105.200 ;
        RECT 43.000 104.200 43.300 104.800 ;
        RECT 40.600 103.800 41.000 104.200 ;
        RECT 43.000 103.800 43.400 104.200 ;
        RECT 48.600 103.200 48.900 104.800 ;
        RECT 49.400 103.200 49.700 105.800 ;
        RECT 51.000 105.100 51.400 105.200 ;
        RECT 51.800 105.100 52.200 105.200 ;
        RECT 51.000 104.800 52.200 105.100 ;
        RECT 50.200 104.100 50.600 104.200 ;
        RECT 51.000 104.100 51.400 104.200 ;
        RECT 50.200 103.800 51.400 104.100 ;
        RECT 48.600 102.800 49.000 103.200 ;
        RECT 49.400 102.800 49.800 103.200 ;
        RECT 51.000 102.800 51.400 103.200 ;
        RECT 47.800 100.800 48.200 101.200 ;
        RECT 45.400 99.800 45.800 100.200 ;
        RECT 45.400 99.200 45.700 99.800 ;
        RECT 47.800 99.200 48.100 100.800 ;
        RECT 51.000 99.200 51.300 102.800 ;
        RECT 45.400 98.800 45.800 99.200 ;
        RECT 47.800 98.800 48.200 99.200 ;
        RECT 51.000 98.800 51.400 99.200 ;
        RECT 40.600 97.800 41.000 98.200 ;
        RECT 46.200 97.800 46.600 98.200 ;
        RECT 50.200 97.800 50.600 98.200 ;
        RECT 40.600 94.200 40.900 97.800 ;
        RECT 44.600 96.800 45.000 97.200 ;
        RECT 41.400 95.100 41.800 95.200 ;
        RECT 42.200 95.100 42.600 95.200 ;
        RECT 41.400 94.800 42.600 95.100 ;
        RECT 44.600 94.200 44.900 96.800 ;
        RECT 46.200 96.200 46.500 97.800 ;
        RECT 48.600 96.800 49.000 97.200 ;
        RECT 46.200 95.800 46.600 96.200 ;
        RECT 47.000 96.100 47.400 96.200 ;
        RECT 47.800 96.100 48.200 96.200 ;
        RECT 47.000 95.800 48.200 96.100 ;
        RECT 45.400 94.800 45.800 95.200 ;
        RECT 47.000 95.100 47.400 95.200 ;
        RECT 47.800 95.100 48.200 95.200 ;
        RECT 47.000 94.800 48.200 95.100 ;
        RECT 40.600 93.800 41.000 94.200 ;
        RECT 42.200 93.800 42.600 94.200 ;
        RECT 44.600 93.800 45.000 94.200 ;
        RECT 45.400 94.100 45.700 94.800 ;
        RECT 46.200 94.100 46.600 94.200 ;
        RECT 45.400 93.800 46.600 94.100 ;
        RECT 40.600 92.200 40.900 93.800 ;
        RECT 40.600 91.800 41.000 92.200 ;
        RECT 42.200 89.200 42.500 93.800 ;
        RECT 43.000 92.800 43.400 93.200 ;
        RECT 45.400 92.800 45.800 93.200 ;
        RECT 43.000 92.200 43.300 92.800 ;
        RECT 43.000 91.800 43.400 92.200 ;
        RECT 45.400 89.200 45.700 92.800 ;
        RECT 42.200 88.800 42.600 89.200 ;
        RECT 45.400 88.800 45.800 89.200 ;
        RECT 47.000 89.100 47.400 89.200 ;
        RECT 47.800 89.100 48.200 89.200 ;
        RECT 47.000 88.800 48.200 89.100 ;
        RECT 43.000 87.100 43.400 87.200 ;
        RECT 43.800 87.100 44.200 87.200 ;
        RECT 43.000 86.800 44.200 87.100 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 44.600 86.200 44.900 86.800 ;
        RECT 40.600 85.800 41.000 86.200 ;
        RECT 43.800 85.800 44.200 86.200 ;
        RECT 44.600 85.800 45.000 86.200 ;
        RECT 40.600 85.200 40.900 85.800 ;
        RECT 40.600 84.800 41.000 85.200 ;
        RECT 39.000 81.800 39.400 82.200 ;
        RECT 39.800 81.800 40.200 82.200 ;
        RECT 39.000 80.200 39.300 81.800 ;
        RECT 39.000 79.800 39.400 80.200 ;
        RECT 35.000 78.800 35.400 79.200 ;
        RECT 31.800 75.100 32.200 75.200 ;
        RECT 31.000 74.800 32.200 75.100 ;
        RECT 23.800 68.800 24.200 69.200 ;
        RECT 27.800 68.800 28.200 69.200 ;
        RECT 28.600 68.800 29.000 69.200 ;
        RECT 27.800 68.200 28.100 68.800 ;
        RECT 28.600 68.200 28.900 68.800 ;
        RECT 25.400 67.800 25.800 68.200 ;
        RECT 26.200 68.100 26.600 68.200 ;
        RECT 27.000 68.100 27.400 68.200 ;
        RECT 26.200 67.800 27.400 68.100 ;
        RECT 27.800 67.800 28.200 68.200 ;
        RECT 28.600 67.800 29.000 68.200 ;
        RECT 25.400 67.200 25.700 67.800 ;
        RECT 19.800 66.800 20.200 67.200 ;
        RECT 22.200 66.800 22.600 67.200 ;
        RECT 23.800 66.800 24.200 67.200 ;
        RECT 25.400 66.800 25.800 67.200 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 27.000 67.100 27.400 67.200 ;
        RECT 26.200 66.800 27.400 67.100 ;
        RECT 19.800 66.200 20.100 66.800 ;
        RECT 22.200 66.200 22.500 66.800 ;
        RECT 23.800 66.200 24.100 66.800 ;
        RECT 19.000 65.800 19.400 66.200 ;
        RECT 19.800 65.800 20.200 66.200 ;
        RECT 21.400 65.800 21.800 66.200 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 23.800 65.800 24.200 66.200 ;
        RECT 19.000 65.200 19.300 65.800 ;
        RECT 19.800 65.200 20.100 65.800 ;
        RECT 19.000 64.800 19.400 65.200 ;
        RECT 19.800 64.800 20.200 65.200 ;
        RECT 19.000 63.800 19.400 64.200 ;
        RECT 16.600 55.100 17.000 55.200 ;
        RECT 13.400 54.700 13.800 55.100 ;
        RECT 15.800 54.800 17.000 55.100 ;
        RECT 13.400 49.200 13.700 54.700 ;
        RECT 16.600 53.200 16.900 54.800 ;
        RECT 16.600 52.800 17.000 53.200 ;
        RECT 17.400 52.100 17.800 57.900 ;
        RECT 17.400 50.800 17.800 51.200 ;
        RECT 13.400 48.800 13.800 49.200 ;
        RECT 17.400 48.200 17.700 50.800 ;
        RECT 19.000 49.200 19.300 63.800 ;
        RECT 21.400 59.200 21.700 65.800 ;
        RECT 23.800 64.800 24.200 65.200 ;
        RECT 23.800 59.200 24.100 64.800 ;
        RECT 20.600 58.800 21.000 59.200 ;
        RECT 21.400 58.800 21.800 59.200 ;
        RECT 23.800 58.800 24.200 59.200 ;
        RECT 20.600 56.200 20.900 58.800 ;
        RECT 22.200 57.100 22.600 57.200 ;
        RECT 23.000 57.100 23.400 57.200 ;
        RECT 22.200 56.800 23.400 57.100 ;
        RECT 27.800 56.800 28.200 57.200 ;
        RECT 27.800 56.200 28.100 56.800 ;
        RECT 20.600 55.800 21.000 56.200 ;
        RECT 24.600 55.800 25.000 56.200 ;
        RECT 27.800 55.800 28.200 56.200 ;
        RECT 22.200 54.800 22.600 55.200 ;
        RECT 22.200 54.200 22.500 54.800 ;
        RECT 24.600 54.200 24.900 55.800 ;
        RECT 28.600 55.200 28.900 67.800 ;
        RECT 30.200 63.100 30.600 68.900 ;
        RECT 31.800 66.200 32.100 74.800 ;
        RECT 32.600 72.100 33.000 77.900 ;
        RECT 39.000 77.800 39.400 78.200 ;
        RECT 37.400 74.800 37.800 75.200 ;
        RECT 37.400 74.200 37.700 74.800 ;
        RECT 37.400 73.800 37.800 74.200 ;
        RECT 39.000 69.200 39.300 77.800 ;
        RECT 31.800 65.800 32.200 66.200 ;
        RECT 32.600 66.100 33.000 66.200 ;
        RECT 33.400 66.100 33.800 66.200 ;
        RECT 32.600 65.800 33.800 66.100 ;
        RECT 25.400 54.800 25.800 55.200 ;
        RECT 26.200 54.800 26.600 55.200 ;
        RECT 28.600 54.800 29.000 55.200 ;
        RECT 30.200 54.800 30.600 55.200 ;
        RECT 22.200 53.800 22.600 54.200 ;
        RECT 24.600 53.800 25.000 54.200 ;
        RECT 21.400 52.800 21.800 53.200 ;
        RECT 19.800 51.800 20.200 52.200 ;
        RECT 20.600 51.800 21.000 52.200 ;
        RECT 19.800 51.200 20.100 51.800 ;
        RECT 19.800 50.800 20.200 51.200 ;
        RECT 19.000 48.800 19.400 49.200 ;
        RECT 10.200 47.800 10.600 48.200 ;
        RECT 16.600 47.800 17.000 48.200 ;
        RECT 17.400 47.800 17.800 48.200 ;
        RECT 8.600 44.800 9.000 45.200 ;
        RECT 9.400 39.100 9.800 39.200 ;
        RECT 10.200 39.100 10.500 47.800 ;
        RECT 16.600 47.200 16.900 47.800 ;
        RECT 12.600 46.800 13.000 47.200 ;
        RECT 16.600 46.800 17.000 47.200 ;
        RECT 17.400 46.800 17.800 47.200 ;
        RECT 12.600 46.200 12.900 46.800 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 15.000 45.800 15.400 46.200 ;
        RECT 15.800 46.100 16.200 46.200 ;
        RECT 16.600 46.100 17.000 46.200 ;
        RECT 15.800 45.800 17.000 46.100 ;
        RECT 15.000 44.200 15.300 45.800 ;
        RECT 15.000 43.800 15.400 44.200 ;
        RECT 9.400 38.800 10.500 39.100 ;
        RECT 11.000 41.800 11.400 42.200 ;
        RECT 3.800 35.800 4.200 36.200 ;
        RECT 3.800 35.100 4.200 35.200 ;
        RECT 4.600 35.100 5.000 35.200 ;
        RECT 3.800 34.800 5.000 35.100 ;
        RECT 3.000 32.800 3.400 33.200 ;
        RECT 0.600 25.100 1.000 27.900 ;
        RECT 2.200 23.100 2.600 28.900 ;
        RECT 3.000 28.200 3.300 32.800 ;
        RECT 7.000 32.100 7.400 37.900 ;
        RECT 11.000 35.200 11.300 41.800 ;
        RECT 14.200 39.800 14.600 40.200 ;
        RECT 13.400 35.800 13.800 36.200 ;
        RECT 13.400 35.200 13.700 35.800 ;
        RECT 14.200 35.200 14.500 39.800 ;
        RECT 17.400 39.200 17.700 46.800 ;
        RECT 19.000 45.100 19.400 45.200 ;
        RECT 19.800 45.100 20.200 45.200 ;
        RECT 19.000 44.800 20.200 45.100 ;
        RECT 20.600 43.200 20.900 51.800 ;
        RECT 21.400 49.200 21.700 52.800 ;
        RECT 21.400 48.800 21.800 49.200 ;
        RECT 23.000 45.800 23.400 46.200 ;
        RECT 20.600 42.800 21.000 43.200 ;
        RECT 20.600 40.200 20.900 42.800 ;
        RECT 20.600 39.800 21.000 40.200 ;
        RECT 17.400 38.800 17.800 39.200 ;
        RECT 18.200 35.800 18.600 36.200 ;
        RECT 18.200 35.200 18.500 35.800 ;
        RECT 10.200 34.800 10.600 35.200 ;
        RECT 11.000 34.800 11.400 35.200 ;
        RECT 13.400 34.800 13.800 35.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 15.000 34.800 15.400 35.200 ;
        RECT 18.200 34.800 18.600 35.200 ;
        RECT 10.200 34.200 10.500 34.800 ;
        RECT 10.200 33.800 10.600 34.200 ;
        RECT 9.400 29.800 9.800 30.200 ;
        RECT 9.400 29.200 9.700 29.800 ;
        RECT 6.200 28.800 6.600 29.200 ;
        RECT 3.000 27.800 3.400 28.200 ;
        RECT 6.200 26.200 6.500 28.800 ;
        RECT 3.800 26.100 4.200 26.200 ;
        RECT 4.600 26.100 5.000 26.200 ;
        RECT 3.800 25.800 5.000 26.100 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 3.800 24.800 4.200 25.200 ;
        RECT 1.400 15.800 1.800 16.200 ;
        RECT 1.400 15.200 1.700 15.800 ;
        RECT 3.800 15.200 4.100 24.800 ;
        RECT 7.000 23.100 7.400 28.900 ;
        RECT 9.400 28.800 9.800 29.200 ;
        RECT 11.800 26.800 12.200 27.200 ;
        RECT 12.600 26.800 13.000 27.200 ;
        RECT 11.800 26.200 12.100 26.800 ;
        RECT 11.800 25.800 12.200 26.200 ;
        RECT 12.600 19.200 12.900 26.800 ;
        RECT 13.400 25.200 13.700 34.800 ;
        RECT 15.000 27.200 15.300 34.800 ;
        RECT 15.800 33.800 16.200 34.200 ;
        RECT 17.400 33.800 17.800 34.200 ;
        RECT 15.800 28.200 16.100 33.800 ;
        RECT 17.400 30.200 17.700 33.800 ;
        RECT 19.000 33.100 19.400 35.900 ;
        RECT 19.000 31.800 19.400 32.200 ;
        RECT 20.600 32.100 21.000 37.900 ;
        RECT 22.200 34.800 22.600 35.200 ;
        RECT 22.200 34.200 22.500 34.800 ;
        RECT 22.200 33.800 22.600 34.200 ;
        RECT 21.400 32.800 21.800 33.200 ;
        RECT 17.400 29.800 17.800 30.200 ;
        RECT 19.000 29.200 19.300 31.800 ;
        RECT 21.400 29.200 21.700 32.800 ;
        RECT 18.200 28.800 18.600 29.200 ;
        RECT 19.000 28.800 19.400 29.200 ;
        RECT 21.400 28.800 21.800 29.200 ;
        RECT 15.800 27.800 16.200 28.200 ;
        RECT 17.400 27.800 17.800 28.200 ;
        RECT 17.400 27.200 17.700 27.800 ;
        RECT 15.000 26.800 15.400 27.200 ;
        RECT 15.800 26.800 16.200 27.200 ;
        RECT 17.400 26.800 17.800 27.200 ;
        RECT 15.800 26.200 16.100 26.800 ;
        RECT 15.000 25.800 15.400 26.200 ;
        RECT 15.800 25.800 16.200 26.200 ;
        RECT 16.600 25.800 17.000 26.200 ;
        RECT 15.000 25.200 15.300 25.800 ;
        RECT 13.400 24.800 13.800 25.200 ;
        RECT 15.000 24.800 15.400 25.200 ;
        RECT 12.600 18.800 13.000 19.200 ;
        RECT 9.400 17.800 9.800 18.200 ;
        RECT 4.600 16.800 5.000 17.200 ;
        RECT 4.600 15.200 4.900 16.800 ;
        RECT 5.400 16.100 5.800 16.200 ;
        RECT 6.200 16.100 6.600 16.200 ;
        RECT 5.400 15.800 6.600 16.100 ;
        RECT 1.400 14.800 1.800 15.200 ;
        RECT 3.800 14.800 4.200 15.200 ;
        RECT 4.600 14.800 5.000 15.200 ;
        RECT 6.200 15.100 6.600 15.200 ;
        RECT 7.000 15.100 7.400 15.200 ;
        RECT 6.200 14.800 7.400 15.100 ;
        RECT 7.800 14.800 8.200 15.200 ;
        RECT 7.800 14.200 8.100 14.800 ;
        RECT 7.800 13.800 8.200 14.200 ;
        RECT 6.200 12.800 6.600 13.200 ;
        RECT 3.000 11.800 3.400 12.200 ;
        RECT 0.600 5.100 1.000 7.900 ;
        RECT 2.200 3.100 2.600 8.900 ;
        RECT 3.000 6.300 3.300 11.800 ;
        RECT 6.200 9.200 6.500 12.800 ;
        RECT 8.600 11.800 9.000 12.200 ;
        RECT 6.200 8.800 6.600 9.200 ;
        RECT 4.600 7.100 5.000 7.200 ;
        RECT 5.400 7.100 5.800 7.200 ;
        RECT 4.600 6.800 5.800 7.100 ;
        RECT 3.000 5.900 3.400 6.300 ;
        RECT 7.000 3.100 7.400 8.900 ;
        RECT 8.600 6.200 8.900 11.800 ;
        RECT 9.400 10.200 9.700 17.800 ;
        RECT 14.200 16.800 14.600 17.200 ;
        RECT 10.200 15.100 10.600 15.200 ;
        RECT 11.000 15.100 11.400 15.200 ;
        RECT 10.200 14.800 11.400 15.100 ;
        RECT 11.800 13.100 12.200 13.200 ;
        RECT 12.600 13.100 13.000 13.200 ;
        RECT 11.800 12.800 13.000 13.100 ;
        RECT 9.400 9.800 9.800 10.200 ;
        RECT 9.400 9.200 9.700 9.800 ;
        RECT 9.400 8.800 9.800 9.200 ;
        RECT 8.600 5.800 9.000 6.200 ;
        RECT 10.200 5.100 10.600 7.900 ;
        RECT 11.000 7.800 11.400 8.200 ;
        RECT 11.000 7.200 11.300 7.800 ;
        RECT 11.000 6.800 11.400 7.200 ;
        RECT 11.800 3.100 12.200 8.900 ;
        RECT 14.200 7.200 14.500 16.800 ;
        RECT 15.000 12.100 15.400 17.900 ;
        RECT 16.600 13.200 16.900 25.800 ;
        RECT 18.200 14.200 18.500 28.800 ;
        RECT 19.000 26.800 19.400 27.200 ;
        RECT 23.000 27.100 23.300 45.800 ;
        RECT 25.400 44.200 25.700 54.800 ;
        RECT 26.200 54.200 26.500 54.800 ;
        RECT 26.200 53.800 26.600 54.200 ;
        RECT 25.400 43.800 25.800 44.200 ;
        RECT 25.400 32.100 25.800 37.900 ;
        RECT 22.200 26.800 23.300 27.100 ;
        RECT 19.000 18.200 19.300 26.800 ;
        RECT 19.800 26.100 20.200 26.200 ;
        RECT 20.600 26.100 21.000 26.200 ;
        RECT 19.800 25.800 21.000 26.100 ;
        RECT 19.000 17.800 19.400 18.200 ;
        RECT 19.000 14.700 19.400 15.100 ;
        RECT 18.200 13.800 18.600 14.200 ;
        RECT 15.800 12.800 16.200 13.200 ;
        RECT 16.600 12.800 17.000 13.200 ;
        RECT 15.800 8.200 16.100 12.800 ;
        RECT 16.600 10.200 16.900 12.800 ;
        RECT 19.000 12.200 19.300 14.700 ;
        RECT 19.000 11.800 19.400 12.200 ;
        RECT 19.800 12.100 20.200 17.900 ;
        RECT 22.200 17.200 22.500 26.800 ;
        RECT 23.000 24.800 23.400 25.200 ;
        RECT 22.200 16.800 22.600 17.200 ;
        RECT 20.600 14.800 21.000 15.200 ;
        RECT 19.800 10.800 20.200 11.200 ;
        RECT 16.600 9.800 17.000 10.200 ;
        RECT 19.000 9.800 19.400 10.200 ;
        RECT 19.000 9.200 19.300 9.800 ;
        RECT 15.800 7.800 16.200 8.200 ;
        RECT 12.600 6.800 13.000 7.200 ;
        RECT 14.200 6.800 14.600 7.200 ;
        RECT 12.600 6.300 12.900 6.800 ;
        RECT 12.600 5.900 13.000 6.300 ;
        RECT 16.600 3.100 17.000 8.900 ;
        RECT 19.000 8.800 19.400 9.200 ;
        RECT 19.800 6.200 20.100 10.800 ;
        RECT 20.600 7.200 20.900 14.800 ;
        RECT 21.400 13.100 21.800 15.900 ;
        RECT 22.200 15.200 22.500 16.800 ;
        RECT 23.000 15.200 23.300 24.800 ;
        RECT 22.200 14.800 22.600 15.200 ;
        RECT 23.000 14.800 23.400 15.200 ;
        RECT 21.400 11.800 21.800 12.200 ;
        RECT 21.400 9.200 21.700 11.800 ;
        RECT 23.000 11.200 23.300 14.800 ;
        RECT 24.600 11.800 25.000 12.200 ;
        RECT 23.000 10.800 23.400 11.200 ;
        RECT 21.400 8.800 21.800 9.200 ;
        RECT 22.200 8.100 22.600 8.200 ;
        RECT 23.000 8.100 23.400 8.200 ;
        RECT 22.200 7.800 23.400 8.100 ;
        RECT 24.600 7.200 24.900 11.800 ;
        RECT 20.600 6.800 21.000 7.200 ;
        RECT 24.600 6.800 25.000 7.200 ;
        RECT 20.600 6.200 20.900 6.800 ;
        RECT 19.800 5.800 20.200 6.200 ;
        RECT 20.600 5.800 21.000 6.200 ;
        RECT 23.800 6.100 24.200 6.200 ;
        RECT 24.600 6.100 25.000 6.200 ;
        RECT 23.800 5.800 25.000 6.100 ;
        RECT 19.800 5.200 20.100 5.800 ;
        RECT 19.800 4.800 20.200 5.200 ;
        RECT 25.400 5.100 25.800 7.900 ;
        RECT 26.200 6.200 26.500 53.800 ;
        RECT 30.200 53.200 30.500 54.800 ;
        RECT 30.200 52.800 30.600 53.200 ;
        RECT 31.000 53.100 31.400 55.900 ;
        RECT 31.800 54.200 32.100 65.800 ;
        RECT 35.000 63.100 35.400 68.900 ;
        RECT 39.000 68.800 39.400 69.200 ;
        RECT 36.600 65.100 37.000 67.900 ;
        RECT 38.200 66.800 38.600 67.200 ;
        RECT 38.200 66.200 38.500 66.800 ;
        RECT 38.200 65.800 38.600 66.200 ;
        RECT 40.600 62.100 40.900 84.800 ;
        RECT 43.000 81.800 43.400 82.200 ;
        RECT 43.000 75.200 43.300 81.800 ;
        RECT 43.800 78.200 44.100 85.800 ;
        RECT 46.200 84.800 46.600 85.200 ;
        RECT 46.200 84.200 46.500 84.800 ;
        RECT 44.600 83.800 45.000 84.200 ;
        RECT 46.200 83.800 46.600 84.200 ;
        RECT 44.600 79.200 44.900 83.800 ;
        RECT 44.600 78.800 45.000 79.200 ;
        RECT 43.800 77.800 44.200 78.200 ;
        RECT 45.400 75.800 45.800 76.200 ;
        RECT 45.400 75.200 45.700 75.800 ;
        RECT 42.200 74.800 42.600 75.200 ;
        RECT 43.000 74.800 43.400 75.200 ;
        RECT 45.400 74.800 45.800 75.200 ;
        RECT 42.200 71.100 42.500 74.800 ;
        RECT 43.800 73.800 44.200 74.200 ;
        RECT 43.800 72.200 44.100 73.800 ;
        RECT 46.200 73.100 46.600 75.900 ;
        RECT 47.000 73.800 47.400 74.200 ;
        RECT 43.800 71.800 44.200 72.200 ;
        RECT 42.200 70.800 43.300 71.100 ;
        RECT 41.400 63.100 41.800 68.900 ;
        RECT 42.200 66.800 42.600 67.200 ;
        RECT 42.200 66.200 42.500 66.800 ;
        RECT 43.000 66.200 43.300 70.800 ;
        RECT 45.400 66.800 45.800 67.200 ;
        RECT 45.400 66.300 45.700 66.800 ;
        RECT 42.200 65.800 42.600 66.200 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 45.400 65.900 45.800 66.300 ;
        RECT 43.800 63.100 44.200 63.200 ;
        RECT 46.200 63.100 46.600 68.900 ;
        RECT 47.000 67.200 47.300 73.800 ;
        RECT 47.800 72.100 48.200 77.900 ;
        RECT 48.600 69.200 48.900 96.800 ;
        RECT 50.200 96.200 50.500 97.800 ;
        RECT 50.200 95.800 50.600 96.200 ;
        RECT 49.400 83.100 49.800 88.900 ;
        RECT 50.200 76.200 50.500 95.800 ;
        RECT 51.800 93.800 52.200 94.200 ;
        RECT 51.800 90.200 52.100 93.800 ;
        RECT 51.800 89.800 52.200 90.200 ;
        RECT 51.800 89.200 52.100 89.800 ;
        RECT 51.800 88.800 52.200 89.200 ;
        RECT 52.600 85.200 52.900 105.800 ;
        RECT 56.600 105.200 56.900 105.800 ;
        RECT 56.600 104.800 57.000 105.200 ;
        RECT 57.400 95.200 57.700 106.800 ;
        RECT 60.600 105.200 60.900 106.800 ;
        RECT 65.400 106.200 65.700 106.800 ;
        RECT 61.400 105.800 61.800 106.200 ;
        RECT 63.000 106.100 63.400 106.200 ;
        RECT 63.800 106.100 64.200 106.200 ;
        RECT 63.000 105.800 64.200 106.100 ;
        RECT 65.400 105.800 65.800 106.200 ;
        RECT 60.600 104.800 61.000 105.200 ;
        RECT 61.400 101.200 61.700 105.800 ;
        RECT 62.200 104.800 62.600 105.200 ;
        RECT 64.600 105.100 65.000 105.200 ;
        RECT 65.400 105.100 65.800 105.200 ;
        RECT 64.600 104.800 65.800 105.100 ;
        RECT 61.400 100.800 61.800 101.200 ;
        RECT 57.400 94.800 57.800 95.200 ;
        RECT 55.800 94.100 56.200 94.200 ;
        RECT 56.600 94.100 57.000 94.200 ;
        RECT 55.800 93.800 57.000 94.100 ;
        RECT 57.400 93.100 57.800 93.200 ;
        RECT 58.200 93.100 58.600 93.200 ;
        RECT 59.000 93.100 59.400 95.900 ;
        RECT 59.800 93.800 60.200 94.200 ;
        RECT 57.400 92.800 58.600 93.100 ;
        RECT 59.800 92.200 60.100 93.800 ;
        RECT 55.000 91.800 55.400 92.200 ;
        RECT 56.600 91.800 57.000 92.200 ;
        RECT 59.800 91.800 60.200 92.200 ;
        RECT 60.600 92.100 61.000 97.900 ;
        RECT 62.200 97.200 62.500 104.800 ;
        RECT 69.400 104.200 69.700 112.800 ;
        RECT 71.000 111.800 71.400 112.200 ;
        RECT 63.800 104.100 64.200 104.200 ;
        RECT 64.600 104.100 65.000 104.200 ;
        RECT 63.800 103.800 65.000 104.100 ;
        RECT 69.400 103.800 69.800 104.200 ;
        RECT 63.000 102.800 63.400 103.200 ;
        RECT 70.200 103.100 70.600 108.900 ;
        RECT 71.000 106.100 71.300 111.800 ;
        RECT 71.800 106.100 72.200 106.200 ;
        RECT 71.000 105.800 72.200 106.100 ;
        RECT 63.000 102.200 63.300 102.800 ;
        RECT 63.000 101.800 63.400 102.200 ;
        RECT 67.800 101.800 68.200 102.200 ;
        RECT 67.800 99.200 68.100 101.800 ;
        RECT 67.800 98.800 68.200 99.200 ;
        RECT 62.200 96.800 62.600 97.200 ;
        RECT 64.600 96.800 65.000 97.200 ;
        RECT 64.600 95.200 64.900 96.800 ;
        RECT 62.200 95.100 62.600 95.200 ;
        RECT 63.000 95.100 63.400 95.200 ;
        RECT 62.200 94.800 63.400 95.100 ;
        RECT 64.600 94.800 65.000 95.200 ;
        RECT 65.400 92.100 65.800 97.900 ;
        RECT 70.200 94.800 70.600 95.200 ;
        RECT 70.200 94.200 70.500 94.800 ;
        RECT 70.200 93.800 70.600 94.200 ;
        RECT 53.400 88.800 53.800 89.200 ;
        RECT 53.400 86.300 53.700 88.800 ;
        RECT 53.400 85.900 53.800 86.300 ;
        RECT 52.600 84.800 53.000 85.200 ;
        RECT 54.200 83.100 54.600 88.900 ;
        RECT 55.000 87.200 55.300 91.800 ;
        RECT 56.600 88.200 56.900 91.800 ;
        RECT 64.600 90.800 65.000 91.200 ;
        RECT 59.800 89.800 60.200 90.200 ;
        RECT 58.200 89.100 58.600 89.200 ;
        RECT 59.000 89.100 59.400 89.200 ;
        RECT 58.200 88.800 59.400 89.100 ;
        RECT 59.800 88.200 60.100 89.800 ;
        RECT 64.600 89.200 64.900 90.800 ;
        RECT 70.200 89.800 70.600 90.200 ;
        RECT 62.200 88.800 62.600 89.200 ;
        RECT 64.600 88.800 65.000 89.200 ;
        RECT 55.000 86.800 55.400 87.200 ;
        RECT 53.400 79.800 53.800 80.200 ;
        RECT 51.800 77.800 52.200 78.200 ;
        RECT 50.200 75.800 50.600 76.200 ;
        RECT 49.400 75.100 49.800 75.200 ;
        RECT 50.200 75.100 50.600 75.200 ;
        RECT 49.400 74.800 50.600 75.100 ;
        RECT 48.600 68.800 49.000 69.200 ;
        RECT 51.800 68.200 52.100 77.800 ;
        RECT 52.600 72.100 53.000 77.900 ;
        RECT 53.400 69.100 53.700 79.800 ;
        RECT 55.000 76.200 55.300 86.800 ;
        RECT 55.800 85.100 56.200 87.900 ;
        RECT 56.600 87.800 57.000 88.200 ;
        RECT 59.800 87.800 60.200 88.200 ;
        RECT 62.200 87.200 62.500 88.800 ;
        RECT 70.200 88.200 70.500 89.800 ;
        RECT 69.400 87.800 69.800 88.200 ;
        RECT 70.200 87.800 70.600 88.200 ;
        RECT 72.600 88.100 72.900 114.800 ;
        RECT 73.400 113.800 73.800 114.200 ;
        RECT 73.400 100.200 73.700 113.800 ;
        RECT 74.200 113.200 74.500 116.800 ;
        RECT 75.000 115.200 75.300 121.800 ;
        RECT 80.600 118.100 80.900 131.800 ;
        RECT 83.800 131.200 84.100 133.800 ;
        RECT 87.800 132.200 88.100 133.800 ;
        RECT 87.800 131.800 88.200 132.200 ;
        RECT 88.600 132.100 89.000 132.200 ;
        RECT 89.400 132.100 89.800 132.200 ;
        RECT 88.600 131.800 89.800 132.100 ;
        RECT 81.400 130.800 81.800 131.200 ;
        RECT 83.800 130.800 84.200 131.200 ;
        RECT 81.400 119.200 81.700 130.800 ;
        RECT 82.200 125.100 82.600 127.900 ;
        RECT 83.800 123.100 84.200 128.900 ;
        RECT 85.400 127.800 85.800 128.200 ;
        RECT 85.400 127.200 85.700 127.800 ;
        RECT 85.400 126.800 85.800 127.200 ;
        RECT 86.200 126.800 86.600 127.200 ;
        RECT 86.200 126.200 86.500 126.800 ;
        RECT 86.200 125.800 86.600 126.200 ;
        RECT 88.600 123.100 89.000 128.900 ;
        RECT 81.400 118.800 81.800 119.200 ;
        RECT 80.600 117.800 81.700 118.100 ;
        RECT 80.600 116.800 81.000 117.200 ;
        RECT 75.000 114.800 75.400 115.200 ;
        RECT 75.800 114.800 76.200 115.200 ;
        RECT 78.200 114.800 78.600 115.200 ;
        RECT 75.800 113.200 76.100 114.800 ;
        RECT 74.200 112.800 74.600 113.200 ;
        RECT 75.800 112.800 76.200 113.200 ;
        RECT 75.000 103.100 75.400 108.900 ;
        RECT 78.200 108.200 78.500 114.800 ;
        RECT 79.000 111.800 79.400 112.200 ;
        RECT 75.800 106.800 76.200 107.200 ;
        RECT 75.800 104.100 76.100 106.800 ;
        RECT 76.600 105.100 77.000 107.900 ;
        RECT 78.200 107.800 78.600 108.200 ;
        RECT 77.400 107.100 77.800 107.200 ;
        RECT 78.200 107.100 78.600 107.200 ;
        RECT 77.400 106.800 78.600 107.100 ;
        RECT 75.800 103.800 76.900 104.100 ;
        RECT 73.400 99.800 73.800 100.200 ;
        RECT 76.600 97.200 76.900 103.800 ;
        RECT 79.000 103.200 79.300 111.800 ;
        RECT 80.600 110.200 80.900 116.800 ;
        RECT 81.400 116.200 81.700 117.800 ;
        RECT 83.000 116.800 83.400 117.200 ;
        RECT 83.000 116.200 83.300 116.800 ;
        RECT 92.600 116.200 92.900 134.800 ;
        RECT 93.400 134.200 93.700 141.800 ;
        RECT 95.800 138.800 96.200 139.200 ;
        RECT 95.800 135.200 96.100 138.800 ;
        RECT 95.800 134.800 96.200 135.200 ;
        RECT 93.400 133.800 93.800 134.200 ;
        RECT 95.000 134.100 95.400 134.200 ;
        RECT 95.800 134.100 96.200 134.200 ;
        RECT 95.000 133.800 96.200 134.100 ;
        RECT 94.200 131.800 94.600 132.200 ;
        RECT 96.600 131.800 97.000 132.200 ;
        RECT 99.000 132.100 99.400 137.900 ;
        RECT 101.400 133.200 101.700 146.800 ;
        RECT 103.800 139.200 104.100 151.800 ;
        RECT 104.600 147.200 104.900 151.800 ;
        RECT 105.400 147.200 105.700 156.800 ;
        RECT 106.200 152.100 106.600 157.900 ;
        RECT 107.000 157.200 107.300 161.800 ;
        RECT 107.000 156.800 107.400 157.200 ;
        RECT 109.400 155.800 109.800 156.200 ;
        RECT 109.400 155.200 109.700 155.800 ;
        RECT 109.400 154.800 109.800 155.200 ;
        RECT 110.200 152.800 110.600 153.200 ;
        RECT 108.600 148.800 109.000 149.200 ;
        RECT 108.600 148.200 108.900 148.800 ;
        RECT 107.000 147.800 107.400 148.200 ;
        RECT 108.600 147.800 109.000 148.200 ;
        RECT 107.000 147.200 107.300 147.800 ;
        RECT 104.600 146.800 105.000 147.200 ;
        RECT 105.400 146.800 105.800 147.200 ;
        RECT 107.000 146.800 107.400 147.200 ;
        RECT 108.600 146.200 108.900 147.800 ;
        RECT 110.200 147.200 110.500 152.800 ;
        RECT 111.000 152.100 111.400 157.900 ;
        RECT 112.600 157.200 112.900 166.800 ;
        RECT 114.200 163.100 114.600 168.900 ;
        RECT 115.800 165.100 116.200 167.900 ;
        RECT 117.400 161.800 117.800 162.200 ;
        RECT 122.200 162.100 122.600 168.900 ;
        RECT 123.000 162.100 123.400 168.900 ;
        RECT 123.800 162.100 124.200 168.900 ;
        RECT 124.600 163.100 125.000 168.900 ;
        RECT 125.400 168.800 125.800 169.200 ;
        RECT 125.400 168.200 125.700 168.800 ;
        RECT 125.400 167.800 125.800 168.200 ;
        RECT 125.400 164.800 125.800 165.200 ;
        RECT 117.400 159.200 117.700 161.800 ;
        RECT 117.400 158.800 117.800 159.200 ;
        RECT 112.600 156.800 113.000 157.200 ;
        RECT 114.200 157.100 114.600 157.200 ;
        RECT 115.000 157.100 115.400 157.200 ;
        RECT 114.200 156.800 115.400 157.100 ;
        RECT 111.800 154.800 112.200 155.200 ;
        RECT 111.800 149.200 112.100 154.800 ;
        RECT 112.600 153.100 113.000 155.900 ;
        RECT 114.200 153.800 114.600 154.200 ;
        RECT 113.400 151.800 113.800 152.200 ;
        RECT 113.400 149.200 113.700 151.800 ;
        RECT 111.800 148.800 112.200 149.200 ;
        RECT 113.400 148.800 113.800 149.200 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 114.200 146.200 114.500 153.800 ;
        RECT 115.800 152.100 116.200 157.900 ;
        RECT 118.200 155.100 118.600 155.200 ;
        RECT 119.000 155.100 119.400 155.200 ;
        RECT 118.200 154.800 119.400 155.100 ;
        RECT 119.000 153.800 119.400 154.200 ;
        RECT 115.000 150.800 115.400 151.200 ;
        RECT 115.000 146.200 115.300 150.800 ;
        RECT 115.800 149.800 116.200 150.200 ;
        RECT 115.800 146.200 116.100 149.800 ;
        RECT 119.000 147.200 119.300 153.800 ;
        RECT 120.600 152.100 121.000 157.900 ;
        RECT 122.200 153.100 122.600 155.900 ;
        RECT 125.400 154.200 125.700 164.800 ;
        RECT 126.200 163.100 126.600 168.900 ;
        RECT 127.000 166.800 127.400 167.200 ;
        RECT 125.400 153.800 125.800 154.200 ;
        RECT 127.000 153.200 127.300 166.800 ;
        RECT 127.800 163.100 128.200 168.900 ;
        RECT 128.600 162.100 129.000 168.900 ;
        RECT 129.400 162.100 129.800 168.900 ;
        RECT 135.800 164.800 136.200 165.200 ;
        RECT 127.800 157.800 128.200 158.200 ;
        RECT 130.200 157.800 130.600 158.200 ;
        RECT 127.800 155.200 128.100 157.800 ;
        RECT 130.200 155.200 130.500 157.800 ;
        RECT 127.800 154.800 128.200 155.200 ;
        RECT 128.600 154.800 129.000 155.200 ;
        RECT 129.400 154.800 129.800 155.200 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 133.400 154.800 133.800 155.200 ;
        RECT 123.000 153.100 123.400 153.200 ;
        RECT 123.800 153.100 124.200 153.200 ;
        RECT 123.000 152.800 124.200 153.100 ;
        RECT 127.000 152.800 127.400 153.200 ;
        RECT 119.000 146.800 119.400 147.200 ;
        RECT 104.600 145.800 105.000 146.200 ;
        RECT 108.600 145.800 109.000 146.200 ;
        RECT 112.600 146.100 113.000 146.200 ;
        RECT 113.400 146.100 113.800 146.200 ;
        RECT 112.600 145.800 113.800 146.100 ;
        RECT 114.200 145.800 114.600 146.200 ;
        RECT 115.000 145.800 115.400 146.200 ;
        RECT 115.800 145.800 116.200 146.200 ;
        RECT 103.800 138.800 104.200 139.200 ;
        RECT 103.000 136.800 103.400 137.200 ;
        RECT 103.000 135.100 103.300 136.800 ;
        RECT 103.000 134.700 103.400 135.100 ;
        RECT 102.200 134.100 102.600 134.200 ;
        RECT 103.000 134.100 103.400 134.200 ;
        RECT 102.200 133.800 103.400 134.100 ;
        RECT 101.400 132.800 101.800 133.200 ;
        RECT 103.800 132.100 104.200 137.900 ;
        RECT 104.600 135.200 104.900 145.800 ;
        RECT 107.000 141.800 107.400 142.200 ;
        RECT 107.000 138.200 107.300 141.800 ;
        RECT 107.000 137.800 107.400 138.200 ;
        RECT 104.600 134.800 105.000 135.200 ;
        RECT 105.400 133.100 105.800 135.900 ;
        RECT 107.800 135.800 108.200 136.200 ;
        RECT 107.800 135.200 108.100 135.800 ;
        RECT 114.200 135.200 114.500 145.800 ;
        RECT 115.000 138.200 115.300 145.800 ;
        RECT 117.400 144.800 117.800 145.200 ;
        RECT 117.400 144.200 117.700 144.800 ;
        RECT 117.400 143.800 117.800 144.200 ;
        RECT 115.000 137.800 115.400 138.200 ;
        RECT 106.200 135.100 106.600 135.200 ;
        RECT 107.000 135.100 107.400 135.200 ;
        RECT 106.200 134.800 107.400 135.100 ;
        RECT 107.800 134.800 108.200 135.200 ;
        RECT 110.200 134.800 110.600 135.200 ;
        RECT 114.200 134.800 114.600 135.200 ;
        RECT 115.000 134.800 115.400 135.200 ;
        RECT 115.800 134.800 116.200 135.200 ;
        RECT 107.000 133.800 107.400 134.200 ;
        RECT 108.600 133.800 109.000 134.200 ;
        RECT 93.400 123.800 93.800 124.200 ;
        RECT 81.400 115.800 81.800 116.200 ;
        RECT 83.000 115.800 83.400 116.200 ;
        RECT 92.600 115.800 93.000 116.200 ;
        RECT 92.600 115.200 92.900 115.800 ;
        RECT 81.400 114.800 81.800 115.200 ;
        RECT 84.600 115.100 85.000 115.200 ;
        RECT 85.400 115.100 85.800 115.200 ;
        RECT 84.600 114.800 85.800 115.100 ;
        RECT 86.200 114.800 86.600 115.200 ;
        RECT 91.000 114.800 91.400 115.200 ;
        RECT 92.600 114.800 93.000 115.200 ;
        RECT 81.400 112.200 81.700 114.800 ;
        RECT 86.200 114.200 86.500 114.800 ;
        RECT 91.000 114.200 91.300 114.800 ;
        RECT 93.400 114.200 93.700 123.800 ;
        RECT 94.200 117.200 94.500 131.800 ;
        RECT 96.600 128.200 96.900 131.800 ;
        RECT 103.800 129.800 104.200 130.200 ;
        RECT 103.800 129.200 104.100 129.800 ;
        RECT 107.000 129.200 107.300 133.800 ;
        RECT 108.600 133.200 108.900 133.800 ;
        RECT 110.200 133.200 110.500 134.800 ;
        RECT 108.600 132.800 109.000 133.200 ;
        RECT 110.200 132.800 110.600 133.200 ;
        RECT 110.200 130.200 110.500 132.800 ;
        RECT 113.400 131.800 113.800 132.200 ;
        RECT 107.800 129.800 108.200 130.200 ;
        RECT 110.200 129.800 110.600 130.200 ;
        RECT 107.800 129.200 108.100 129.800 ;
        RECT 103.800 128.800 104.200 129.200 ;
        RECT 107.000 128.800 107.400 129.200 ;
        RECT 107.800 128.800 108.200 129.200 ;
        RECT 96.600 127.800 97.000 128.200 ;
        RECT 106.200 128.100 106.600 128.200 ;
        RECT 107.000 128.100 107.400 128.200 ;
        RECT 106.200 127.800 107.400 128.100 ;
        RECT 95.000 127.100 95.400 127.200 ;
        RECT 95.800 127.100 96.200 127.200 ;
        RECT 95.000 126.800 96.200 127.100 ;
        RECT 96.600 121.200 96.900 127.800 ;
        RECT 99.800 126.800 100.200 127.200 ;
        RECT 101.400 127.100 101.800 127.200 ;
        RECT 102.200 127.100 102.600 127.200 ;
        RECT 101.400 126.800 102.600 127.100 ;
        RECT 103.000 126.800 103.400 127.200 ;
        RECT 99.800 126.200 100.100 126.800 ;
        RECT 103.000 126.200 103.300 126.800 ;
        RECT 98.200 125.800 98.600 126.200 ;
        RECT 99.000 125.800 99.400 126.200 ;
        RECT 99.800 125.800 100.200 126.200 ;
        RECT 102.200 125.800 102.600 126.200 ;
        RECT 103.000 125.800 103.400 126.200 ;
        RECT 105.400 126.100 105.800 126.200 ;
        RECT 106.200 126.100 106.600 126.200 ;
        RECT 105.400 125.800 106.600 126.100 ;
        RECT 96.600 120.800 97.000 121.200 ;
        RECT 95.800 118.800 96.200 119.200 ;
        RECT 95.800 118.200 96.100 118.800 ;
        RECT 95.800 117.800 96.200 118.200 ;
        RECT 97.400 117.800 97.800 118.200 ;
        RECT 94.200 116.800 94.600 117.200 ;
        RECT 95.800 116.800 96.200 117.200 ;
        RECT 96.600 116.800 97.000 117.200 ;
        RECT 95.800 114.200 96.100 116.800 ;
        RECT 96.600 115.200 96.900 116.800 ;
        RECT 97.400 116.200 97.700 117.800 ;
        RECT 97.400 115.800 97.800 116.200 ;
        RECT 96.600 114.800 97.000 115.200 ;
        RECT 83.000 113.800 83.400 114.200 ;
        RECT 84.600 114.100 85.000 114.200 ;
        RECT 84.600 113.800 85.700 114.100 ;
        RECT 86.200 113.800 86.600 114.200 ;
        RECT 91.000 113.800 91.400 114.200 ;
        RECT 93.400 113.800 93.800 114.200 ;
        RECT 95.800 113.800 96.200 114.200 ;
        RECT 83.000 113.200 83.300 113.800 ;
        RECT 83.000 112.800 83.400 113.200 ;
        RECT 81.400 111.800 81.800 112.200 ;
        RECT 80.600 109.800 81.000 110.200 ;
        RECT 85.400 109.200 85.700 113.800 ;
        RECT 92.600 113.100 93.000 113.200 ;
        RECT 93.400 113.100 93.800 113.200 ;
        RECT 92.600 112.800 93.800 113.100 ;
        RECT 87.800 111.800 88.200 112.200 ;
        RECT 87.800 109.200 88.100 111.800 ;
        RECT 85.400 108.800 85.800 109.200 ;
        RECT 87.800 108.800 88.200 109.200 ;
        RECT 82.200 107.800 82.600 108.200 ;
        RECT 82.200 107.200 82.500 107.800 ;
        RECT 82.200 106.800 82.600 107.200 ;
        RECT 83.000 106.800 83.400 107.200 ;
        RECT 86.200 106.800 86.600 107.200 ;
        RECT 91.000 106.800 91.400 107.200 ;
        RECT 79.800 105.800 80.200 106.200 ;
        RECT 82.200 105.800 82.600 106.200 ;
        RECT 79.000 102.800 79.400 103.200 ;
        RECT 76.600 96.800 77.000 97.200 ;
        RECT 73.400 95.800 73.800 96.200 ;
        RECT 73.400 95.200 73.700 95.800 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 73.400 93.800 73.800 94.200 ;
        RECT 73.400 89.200 73.700 93.800 ;
        RECT 74.200 92.200 74.500 94.800 ;
        RECT 74.200 91.800 74.600 92.200 ;
        RECT 75.000 91.800 75.400 92.200 ;
        RECT 75.800 91.800 76.200 92.200 ;
        RECT 77.400 92.100 77.800 97.900 ;
        RECT 75.000 90.200 75.300 91.800 ;
        RECT 75.000 89.800 75.400 90.200 ;
        RECT 73.400 88.800 73.800 89.200 ;
        RECT 72.600 87.800 73.700 88.100 ;
        RECT 69.400 87.200 69.700 87.800 ;
        RECT 56.600 86.800 57.000 87.200 ;
        RECT 57.400 86.800 57.800 87.200 ;
        RECT 62.200 86.800 62.600 87.200 ;
        RECT 66.200 86.800 66.600 87.200 ;
        RECT 67.800 87.100 68.200 87.200 ;
        RECT 68.600 87.100 69.000 87.200 ;
        RECT 67.800 86.800 69.000 87.100 ;
        RECT 69.400 86.800 69.800 87.200 ;
        RECT 56.600 86.200 56.900 86.800 ;
        RECT 57.400 86.200 57.700 86.800 ;
        RECT 66.200 86.200 66.500 86.800 ;
        RECT 70.200 86.200 70.500 87.800 ;
        RECT 56.600 85.800 57.000 86.200 ;
        RECT 57.400 85.800 57.800 86.200 ;
        RECT 61.400 86.100 61.800 86.200 ;
        RECT 62.200 86.100 62.600 86.200 ;
        RECT 61.400 85.800 62.600 86.100 ;
        RECT 66.200 85.800 66.600 86.200 ;
        RECT 67.800 85.800 68.200 86.200 ;
        RECT 70.200 85.800 70.600 86.200 ;
        RECT 71.800 85.800 72.200 86.200 ;
        RECT 56.600 83.200 56.900 85.800 ;
        RECT 56.600 82.800 57.000 83.200 ;
        RECT 55.800 76.800 56.200 77.200 ;
        RECT 57.400 76.800 57.800 77.200 ;
        RECT 55.800 76.200 56.100 76.800 ;
        RECT 55.000 75.800 55.400 76.200 ;
        RECT 55.800 75.800 56.200 76.200 ;
        RECT 57.400 74.200 57.700 76.800 ;
        RECT 57.400 73.800 57.800 74.200 ;
        RECT 54.200 72.100 54.600 72.200 ;
        RECT 55.000 72.100 55.400 72.200 ;
        RECT 54.200 71.800 55.400 72.100 ;
        RECT 55.800 71.800 56.200 72.200 ;
        RECT 59.800 71.800 60.200 72.200 ;
        RECT 60.600 72.100 61.000 77.900 ;
        RECT 61.400 75.800 61.800 76.200 ;
        RECT 61.400 75.200 61.700 75.800 ;
        RECT 61.400 74.800 61.800 75.200 ;
        RECT 55.800 70.200 56.100 71.800 ;
        RECT 57.400 70.800 57.800 71.200 ;
        RECT 55.800 69.800 56.200 70.200 ;
        RECT 53.400 68.800 54.500 69.100 ;
        RECT 47.000 66.800 47.400 67.200 ;
        RECT 47.800 65.100 48.200 67.900 ;
        RECT 48.600 67.800 49.000 68.200 ;
        RECT 51.800 67.800 52.200 68.200 ;
        RECT 53.400 67.800 53.800 68.200 ;
        RECT 48.600 67.200 48.900 67.800 ;
        RECT 48.600 66.800 49.000 67.200 ;
        RECT 50.200 67.100 50.600 67.200 ;
        RECT 51.000 67.100 51.400 67.200 ;
        RECT 50.200 66.800 51.400 67.100 ;
        RECT 53.400 66.200 53.700 67.800 ;
        RECT 54.200 67.200 54.500 68.800 ;
        RECT 55.000 67.800 55.400 68.200 ;
        RECT 55.000 67.200 55.300 67.800 ;
        RECT 54.200 66.800 54.600 67.200 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 48.600 66.100 49.000 66.200 ;
        RECT 49.400 66.100 49.800 66.200 ;
        RECT 48.600 65.800 49.800 66.100 ;
        RECT 53.400 65.800 53.800 66.200 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 56.600 64.200 56.900 65.800 ;
        RECT 56.600 63.800 57.000 64.200 ;
        RECT 43.000 62.800 44.200 63.100 ;
        RECT 47.800 62.800 48.200 63.200 ;
        RECT 40.600 61.800 41.700 62.100 ;
        RECT 31.800 53.800 32.200 54.200 ;
        RECT 31.800 53.200 32.100 53.800 ;
        RECT 31.800 52.800 32.200 53.200 ;
        RECT 32.600 52.100 33.000 57.900 ;
        RECT 33.400 55.800 33.800 56.200 ;
        RECT 33.400 55.100 33.700 55.800 ;
        RECT 33.400 54.700 33.800 55.100 ;
        RECT 36.600 53.800 37.000 54.200 ;
        RECT 35.000 48.800 35.400 49.200 ;
        RECT 35.000 48.200 35.300 48.800 ;
        RECT 35.000 47.800 35.400 48.200 ;
        RECT 27.800 46.800 28.200 47.200 ;
        RECT 31.800 46.800 32.200 47.200 ;
        RECT 27.800 46.200 28.100 46.800 ;
        RECT 31.800 46.200 32.100 46.800 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 28.600 45.800 29.000 46.200 ;
        RECT 31.800 45.800 32.200 46.200 ;
        RECT 28.600 42.200 28.900 45.800 ;
        RECT 35.800 45.100 36.200 47.900 ;
        RECT 36.600 47.200 36.900 53.800 ;
        RECT 37.400 52.100 37.800 57.900 ;
        RECT 40.600 56.800 41.000 57.200 ;
        RECT 40.600 55.200 40.900 56.800 ;
        RECT 40.600 54.800 41.000 55.200 ;
        RECT 41.400 50.200 41.700 61.800 ;
        RECT 43.000 54.200 43.300 62.800 ;
        RECT 47.800 59.200 48.100 62.800 ;
        RECT 52.600 59.800 53.000 60.200 ;
        RECT 52.600 59.200 52.900 59.800 ;
        RECT 47.800 58.800 48.200 59.200 ;
        RECT 52.600 58.800 53.000 59.200 ;
        RECT 44.600 57.800 45.000 58.200 ;
        RECT 44.600 57.200 44.900 57.800 ;
        RECT 44.600 56.800 45.000 57.200 ;
        RECT 46.200 57.100 46.600 57.200 ;
        RECT 47.000 57.100 47.400 57.200 ;
        RECT 46.200 56.800 47.400 57.100 ;
        RECT 56.600 56.800 57.000 57.200 ;
        RECT 48.600 55.800 49.000 56.200 ;
        RECT 49.400 56.100 49.800 56.200 ;
        RECT 50.200 56.100 50.600 56.200 ;
        RECT 49.400 55.800 50.600 56.100 ;
        RECT 55.800 55.800 56.200 56.200 ;
        RECT 45.400 54.800 45.800 55.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 47.800 55.100 48.200 55.200 ;
        RECT 47.000 54.800 48.200 55.100 ;
        RECT 43.000 53.800 43.400 54.200 ;
        RECT 44.600 53.800 45.000 54.200 ;
        RECT 41.400 49.800 41.800 50.200 ;
        RECT 36.600 46.800 37.000 47.200 ;
        RECT 35.800 43.800 36.200 44.200 ;
        RECT 28.600 41.800 29.000 42.200 ;
        RECT 27.800 37.100 28.200 37.200 ;
        RECT 28.600 37.100 29.000 37.200 ;
        RECT 27.800 36.800 29.000 37.100 ;
        RECT 34.200 36.800 34.600 37.200 ;
        RECT 28.600 35.800 29.000 36.200 ;
        RECT 28.600 35.200 28.900 35.800 ;
        RECT 28.600 34.800 29.000 35.200 ;
        RECT 29.400 34.800 29.800 35.200 ;
        RECT 29.400 33.200 29.700 34.800 ;
        RECT 30.200 33.800 30.600 34.200 ;
        RECT 30.200 33.200 30.500 33.800 ;
        RECT 34.200 33.200 34.500 36.800 ;
        RECT 35.000 35.800 35.400 36.200 ;
        RECT 35.000 35.200 35.300 35.800 ;
        RECT 35.800 35.200 36.100 43.800 ;
        RECT 37.400 43.100 37.800 48.900 ;
        RECT 38.200 46.800 38.600 47.200 ;
        RECT 38.200 46.300 38.500 46.800 ;
        RECT 38.200 45.900 38.600 46.300 ;
        RECT 40.600 35.800 41.000 36.200 ;
        RECT 35.000 34.800 35.400 35.200 ;
        RECT 35.800 34.800 36.200 35.200 ;
        RECT 29.400 32.800 29.800 33.200 ;
        RECT 30.200 32.800 30.600 33.200 ;
        RECT 34.200 32.800 34.600 33.200 ;
        RECT 36.600 32.800 37.000 33.200 ;
        RECT 36.600 29.200 36.900 32.800 ;
        RECT 37.400 31.800 37.800 32.200 ;
        RECT 37.400 29.200 37.700 31.800 ;
        RECT 40.600 29.200 40.900 35.800 ;
        RECT 28.600 28.800 29.000 29.200 ;
        RECT 27.800 25.100 28.200 27.900 ;
        RECT 28.600 27.200 28.900 28.800 ;
        RECT 28.600 26.800 29.000 27.200 ;
        RECT 29.400 23.100 29.800 28.900 ;
        RECT 31.000 28.800 31.400 29.200 ;
        RECT 31.000 26.200 31.300 28.800 ;
        RECT 31.000 25.800 31.400 26.200 ;
        RECT 33.400 25.800 33.800 26.200 ;
        RECT 27.800 12.800 28.200 13.200 ;
        RECT 28.600 13.100 29.000 15.900 ;
        RECT 29.400 13.800 29.800 14.200 ;
        RECT 27.800 9.200 28.100 12.800 ;
        RECT 26.200 5.800 26.600 6.200 ;
        RECT 27.000 3.100 27.400 8.900 ;
        RECT 27.800 8.800 28.200 9.200 ;
        RECT 29.400 7.200 29.700 13.800 ;
        RECT 30.200 12.100 30.600 17.900 ;
        RECT 33.400 15.200 33.700 25.800 ;
        RECT 34.200 23.100 34.600 28.900 ;
        RECT 36.600 28.800 37.000 29.200 ;
        RECT 37.400 28.800 37.800 29.200 ;
        RECT 40.600 28.800 41.000 29.200 ;
        RECT 41.400 28.100 41.700 49.800 ;
        RECT 42.200 43.100 42.600 48.900 ;
        RECT 42.200 33.800 42.600 34.200 ;
        RECT 42.200 33.200 42.500 33.800 ;
        RECT 42.200 32.800 42.600 33.200 ;
        RECT 40.600 27.800 41.700 28.100 ;
        RECT 43.000 28.200 43.300 53.800 ;
        RECT 44.600 51.200 44.900 53.800 ;
        RECT 44.600 50.800 45.000 51.200 ;
        RECT 45.400 50.200 45.700 54.800 ;
        RECT 48.600 53.200 48.900 55.800 ;
        RECT 55.800 55.200 56.100 55.800 ;
        RECT 56.600 55.200 56.900 56.800 ;
        RECT 49.400 54.800 49.800 55.200 ;
        RECT 51.800 54.800 52.200 55.200 ;
        RECT 54.200 54.800 54.600 55.200 ;
        RECT 55.800 54.800 56.200 55.200 ;
        RECT 56.600 54.800 57.000 55.200 ;
        RECT 49.400 54.200 49.700 54.800 ;
        RECT 51.800 54.200 52.100 54.800 ;
        RECT 49.400 53.800 49.800 54.200 ;
        RECT 51.800 53.800 52.200 54.200 ;
        RECT 53.400 54.100 53.800 54.200 ;
        RECT 52.600 53.800 53.800 54.100 ;
        RECT 48.600 52.800 49.000 53.200 ;
        RECT 50.200 52.800 50.600 53.200 ;
        RECT 51.000 52.800 51.400 53.200 ;
        RECT 45.400 49.800 45.800 50.200 ;
        RECT 43.800 49.100 44.200 49.200 ;
        RECT 44.600 49.100 45.000 49.200 ;
        RECT 43.800 48.800 45.000 49.100 ;
        RECT 44.600 39.800 45.000 40.200 ;
        RECT 44.600 39.200 44.900 39.800 ;
        RECT 50.200 39.200 50.500 52.800 ;
        RECT 51.000 49.200 51.300 52.800 ;
        RECT 51.000 48.800 51.400 49.200 ;
        RECT 52.600 48.200 52.900 53.800 ;
        RECT 54.200 53.200 54.500 54.800 ;
        RECT 54.200 52.800 54.600 53.200 ;
        RECT 55.000 51.800 55.400 52.200 ;
        RECT 55.800 51.800 56.200 52.200 ;
        RECT 53.400 49.800 53.800 50.200 ;
        RECT 53.400 49.200 53.700 49.800 ;
        RECT 53.400 48.800 53.800 49.200 ;
        RECT 55.000 48.200 55.300 51.800 ;
        RECT 55.800 49.200 56.100 51.800 ;
        RECT 55.800 48.800 56.200 49.200 ;
        RECT 52.600 47.800 53.000 48.200 ;
        RECT 55.000 47.800 55.400 48.200 ;
        RECT 52.600 47.200 52.900 47.800 ;
        RECT 52.600 46.800 53.000 47.200 ;
        RECT 55.000 46.800 55.400 47.200 ;
        RECT 56.600 46.800 57.000 47.200 ;
        RECT 54.200 46.100 54.600 46.200 ;
        RECT 53.400 45.800 54.600 46.100 ;
        RECT 44.600 38.800 45.000 39.200 ;
        RECT 50.200 38.800 50.600 39.200 ;
        RECT 43.800 36.800 44.200 37.200 ;
        RECT 46.200 36.800 46.600 37.200 ;
        RECT 47.800 37.100 48.200 37.200 ;
        RECT 48.600 37.100 49.000 37.200 ;
        RECT 47.800 36.800 49.000 37.100 ;
        RECT 51.000 36.800 51.400 37.200 ;
        RECT 43.800 32.200 44.100 36.800 ;
        RECT 46.200 36.200 46.500 36.800 ;
        RECT 46.200 35.800 46.600 36.200 ;
        RECT 44.600 35.100 45.000 35.200 ;
        RECT 44.600 34.800 45.700 35.100 ;
        RECT 43.800 31.800 44.200 32.200 ;
        RECT 45.400 29.200 45.700 34.800 ;
        RECT 47.000 34.800 47.400 35.200 ;
        RECT 49.400 34.800 49.800 35.200 ;
        RECT 50.200 34.800 50.600 35.200 ;
        RECT 47.000 34.200 47.300 34.800 ;
        RECT 47.000 33.800 47.400 34.200 ;
        RECT 49.400 33.200 49.700 34.800 ;
        RECT 50.200 34.200 50.500 34.800 ;
        RECT 50.200 33.800 50.600 34.200 ;
        RECT 49.400 32.800 49.800 33.200 ;
        RECT 45.400 28.800 45.800 29.200 ;
        RECT 43.000 27.800 43.400 28.200 ;
        RECT 37.400 26.800 37.800 27.200 ;
        RECT 37.400 22.200 37.700 26.800 ;
        RECT 40.600 26.200 40.900 27.800 ;
        RECT 43.000 27.200 43.300 27.800 ;
        RECT 41.400 26.800 41.800 27.200 ;
        RECT 43.000 26.800 43.400 27.200 ;
        RECT 44.600 27.100 45.000 27.200 ;
        RECT 45.400 27.100 45.800 27.200 ;
        RECT 44.600 26.800 45.800 27.100 ;
        RECT 47.000 26.800 47.400 27.200 ;
        RECT 40.600 25.800 41.000 26.200 ;
        RECT 34.200 21.800 34.600 22.200 ;
        RECT 37.400 21.800 37.800 22.200 ;
        RECT 31.800 14.800 32.200 15.200 ;
        RECT 33.400 14.800 33.800 15.200 ;
        RECT 31.800 14.200 32.100 14.800 ;
        RECT 31.800 13.800 32.200 14.200 ;
        RECT 34.200 9.200 34.500 21.800 ;
        RECT 41.400 19.200 41.700 26.800 ;
        RECT 44.600 25.800 45.000 26.200 ;
        RECT 42.200 24.800 42.600 25.200 ;
        RECT 42.200 24.200 42.500 24.800 ;
        RECT 42.200 23.800 42.600 24.200 ;
        RECT 37.400 18.800 37.800 19.200 ;
        RECT 41.400 18.800 41.800 19.200 ;
        RECT 35.000 12.100 35.400 17.900 ;
        RECT 37.400 17.200 37.700 18.800 ;
        RECT 37.400 16.800 37.800 17.200 ;
        RECT 37.400 13.200 37.700 16.800 ;
        RECT 39.000 15.100 39.400 15.200 ;
        RECT 39.800 15.100 40.200 15.200 ;
        RECT 39.000 14.800 40.200 15.100 ;
        RECT 40.600 15.100 41.000 15.200 ;
        RECT 41.400 15.100 41.800 15.200 ;
        RECT 40.600 14.800 41.800 15.100 ;
        RECT 44.600 15.100 44.900 25.800 ;
        RECT 45.400 25.100 45.800 25.200 ;
        RECT 46.200 25.100 46.600 25.200 ;
        RECT 45.400 24.800 46.600 25.100 ;
        RECT 46.200 19.100 46.600 19.200 ;
        RECT 47.000 19.100 47.300 26.800 ;
        RECT 48.600 25.800 49.000 26.200 ;
        RECT 49.400 26.100 49.800 26.200 ;
        RECT 50.200 26.100 50.500 33.800 ;
        RECT 49.400 25.800 50.500 26.100 ;
        RECT 51.000 26.200 51.300 36.800 ;
        RECT 53.400 34.200 53.700 45.800 ;
        RECT 55.000 39.200 55.300 46.800 ;
        RECT 55.000 38.800 55.400 39.200 ;
        RECT 54.200 36.800 54.600 37.200 ;
        RECT 55.000 37.100 55.400 37.200 ;
        RECT 55.800 37.100 56.200 37.200 ;
        RECT 55.000 36.800 56.200 37.100 ;
        RECT 54.200 36.200 54.500 36.800 ;
        RECT 54.200 35.800 54.600 36.200 ;
        RECT 55.000 35.800 55.400 36.200 ;
        RECT 55.000 35.200 55.300 35.800 ;
        RECT 55.000 34.800 55.400 35.200 ;
        RECT 52.600 33.800 53.000 34.200 ;
        RECT 53.400 33.800 53.800 34.200 ;
        RECT 52.600 33.200 52.900 33.800 ;
        RECT 53.400 33.200 53.700 33.800 ;
        RECT 52.600 32.800 53.000 33.200 ;
        RECT 53.400 32.800 53.800 33.200 ;
        RECT 53.400 31.800 53.800 32.200 ;
        RECT 53.400 29.200 53.700 31.800 ;
        RECT 53.400 28.800 53.800 29.200 ;
        RECT 55.000 28.800 55.400 29.200 ;
        RECT 55.000 26.200 55.300 28.800 ;
        RECT 51.000 25.800 51.400 26.200 ;
        RECT 51.800 25.800 52.200 26.200 ;
        RECT 54.200 26.100 54.600 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 54.200 25.800 55.400 26.100 ;
        RECT 48.600 24.200 48.900 25.800 ;
        RECT 50.200 24.800 50.600 25.200 ;
        RECT 51.000 24.800 51.400 25.200 ;
        RECT 48.600 23.800 49.000 24.200 ;
        RECT 49.400 23.800 49.800 24.200 ;
        RECT 49.400 23.200 49.700 23.800 ;
        RECT 50.200 23.200 50.500 24.800 ;
        RECT 49.400 22.800 49.800 23.200 ;
        RECT 50.200 22.800 50.600 23.200 ;
        RECT 51.000 22.200 51.300 24.800 ;
        RECT 51.800 22.200 52.100 25.800 ;
        RECT 49.400 22.100 49.800 22.200 ;
        RECT 50.200 22.100 50.600 22.200 ;
        RECT 49.400 21.800 50.600 22.100 ;
        RECT 51.000 21.800 51.400 22.200 ;
        RECT 51.800 21.800 52.200 22.200 ;
        RECT 46.200 18.800 47.300 19.100 ;
        RECT 44.600 14.800 45.700 15.100 ;
        RECT 41.400 13.800 41.800 14.200 ;
        RECT 44.600 13.800 45.000 14.200 ;
        RECT 41.400 13.200 41.700 13.800 ;
        RECT 44.600 13.200 44.900 13.800 ;
        RECT 37.400 12.800 37.800 13.200 ;
        RECT 41.400 12.800 41.800 13.200 ;
        RECT 44.600 12.800 45.000 13.200 ;
        RECT 45.400 9.200 45.700 14.800 ;
        RECT 48.600 12.100 49.000 17.900 ;
        RECT 51.000 14.800 51.400 15.200 ;
        RECT 49.400 13.800 49.800 14.200 ;
        RECT 49.400 13.200 49.700 13.800 ;
        RECT 49.400 12.800 49.800 13.200 ;
        RECT 33.400 9.100 33.800 9.200 ;
        RECT 34.200 9.100 34.600 9.200 ;
        RECT 27.800 6.800 28.200 7.200 ;
        RECT 29.400 6.800 29.800 7.200 ;
        RECT 27.800 6.300 28.100 6.800 ;
        RECT 27.800 5.900 28.200 6.300 ;
        RECT 31.800 3.100 32.200 8.900 ;
        RECT 33.400 8.800 34.600 9.100 ;
        RECT 36.600 5.100 37.000 7.900 ;
        RECT 37.400 7.800 37.800 8.200 ;
        RECT 37.400 7.200 37.700 7.800 ;
        RECT 37.400 6.800 37.800 7.200 ;
        RECT 38.200 3.100 38.600 8.900 ;
        RECT 41.400 7.800 41.800 8.200 ;
        RECT 41.400 6.200 41.700 7.800 ;
        RECT 41.400 5.800 41.800 6.200 ;
        RECT 43.000 3.100 43.400 8.900 ;
        RECT 45.400 8.800 45.800 9.200 ;
        RECT 49.400 8.800 49.800 9.200 ;
        RECT 49.400 8.200 49.700 8.800 ;
        RECT 49.400 7.800 49.800 8.200 ;
        RECT 50.200 6.800 50.600 7.200 ;
        RECT 50.200 6.200 50.500 6.800 ;
        RECT 51.000 6.200 51.300 14.800 ;
        RECT 52.600 14.700 53.000 15.100 ;
        RECT 52.600 14.200 52.900 14.700 ;
        RECT 52.600 13.800 53.000 14.200 ;
        RECT 52.600 12.800 53.000 13.200 ;
        RECT 52.600 8.200 52.900 12.800 ;
        RECT 53.400 12.100 53.800 17.900 ;
        RECT 55.000 13.100 55.400 15.900 ;
        RECT 56.600 15.100 56.900 46.800 ;
        RECT 57.400 46.200 57.700 70.800 ;
        RECT 59.800 68.200 60.100 71.800 ;
        RECT 59.800 67.800 60.200 68.200 ;
        RECT 62.200 67.200 62.500 85.800 ;
        RECT 63.800 85.100 64.200 85.200 ;
        RECT 64.600 85.100 65.000 85.200 ;
        RECT 63.800 84.800 65.000 85.100 ;
        RECT 64.600 84.100 65.000 84.200 ;
        RECT 65.400 84.100 65.800 84.200 ;
        RECT 64.600 83.800 65.800 84.100 ;
        RECT 66.200 82.200 66.500 85.800 ;
        RECT 67.800 85.200 68.100 85.800 ;
        RECT 67.800 84.800 68.200 85.200 ;
        RECT 69.400 84.800 69.800 85.200 ;
        RECT 69.400 84.200 69.700 84.800 ;
        RECT 69.400 83.800 69.800 84.200 ;
        RECT 71.800 82.200 72.100 85.800 ;
        RECT 63.000 81.800 63.400 82.200 ;
        RECT 66.200 81.800 66.600 82.200 ;
        RECT 69.400 81.800 69.800 82.200 ;
        RECT 71.800 81.800 72.200 82.200 ;
        RECT 63.000 78.200 63.300 81.800 ;
        RECT 63.000 77.800 63.400 78.200 ;
        RECT 63.000 74.800 63.400 75.200 ;
        RECT 63.800 74.800 64.200 75.200 ;
        RECT 63.000 73.200 63.300 74.800 ;
        RECT 63.000 72.800 63.400 73.200 ;
        RECT 63.800 69.200 64.100 74.800 ;
        RECT 64.600 72.800 65.000 73.200 ;
        RECT 64.600 70.200 64.900 72.800 ;
        RECT 65.400 72.100 65.800 77.900 ;
        RECT 66.200 75.800 66.600 76.200 ;
        RECT 64.600 69.800 65.000 70.200 ;
        RECT 63.800 68.800 64.200 69.200 ;
        RECT 62.200 66.800 62.600 67.200 ;
        RECT 63.800 67.100 64.200 67.200 ;
        RECT 64.600 67.100 65.000 67.200 ;
        RECT 63.800 66.800 65.000 67.100 ;
        RECT 62.200 66.200 62.500 66.800 ;
        RECT 66.200 66.200 66.500 75.800 ;
        RECT 67.000 73.100 67.400 75.900 ;
        RECT 69.400 75.200 69.700 81.800 ;
        RECT 72.600 79.800 73.000 80.200 ;
        RECT 72.600 75.200 72.900 79.800 ;
        RECT 73.400 78.200 73.700 87.800 ;
        RECT 74.200 86.800 74.600 87.200 ;
        RECT 74.200 82.200 74.500 86.800 ;
        RECT 75.800 86.200 76.100 91.800 ;
        RECT 79.800 87.200 80.100 105.800 ;
        RECT 82.200 99.100 82.500 105.800 ;
        RECT 83.000 102.200 83.300 106.800 ;
        RECT 83.000 101.800 83.400 102.200 ;
        RECT 86.200 100.200 86.500 106.800 ;
        RECT 87.000 105.800 87.400 106.200 ;
        RECT 86.200 99.800 86.600 100.200 ;
        RECT 81.400 98.800 82.500 99.100 ;
        RECT 86.200 99.100 86.600 99.200 ;
        RECT 87.000 99.100 87.300 105.800 ;
        RECT 86.200 98.800 87.300 99.100 ;
        RECT 87.800 104.800 88.200 105.200 ;
        RECT 81.400 97.200 81.700 98.800 ;
        RECT 87.800 98.200 88.100 104.800 ;
        RECT 91.000 99.200 91.300 106.800 ;
        RECT 92.600 101.800 93.000 102.200 ;
        RECT 91.000 98.800 91.400 99.200 ;
        RECT 81.400 96.800 81.800 97.200 ;
        RECT 80.600 94.800 81.000 95.200 ;
        RECT 80.600 94.200 80.900 94.800 ;
        RECT 80.600 93.800 81.000 94.200 ;
        RECT 79.800 86.800 80.200 87.200 ;
        RECT 75.000 85.800 75.400 86.200 ;
        RECT 75.800 85.800 76.200 86.200 ;
        RECT 76.600 86.100 77.000 86.200 ;
        RECT 77.400 86.100 77.800 86.200 ;
        RECT 76.600 85.800 77.800 86.100 ;
        RECT 79.000 85.800 79.400 86.200 ;
        RECT 75.000 83.100 75.300 85.800 ;
        RECT 76.600 83.800 77.000 84.200 ;
        RECT 75.000 82.800 76.100 83.100 ;
        RECT 74.200 81.800 74.600 82.200 ;
        RECT 75.800 81.200 76.100 82.800 ;
        RECT 75.800 80.800 76.200 81.200 ;
        RECT 74.200 78.800 74.600 79.200 ;
        RECT 74.200 78.200 74.500 78.800 ;
        RECT 73.400 77.800 73.800 78.200 ;
        RECT 74.200 77.800 74.600 78.200 ;
        RECT 73.400 77.200 73.700 77.800 ;
        RECT 76.600 77.200 76.900 83.800 ;
        RECT 73.400 76.800 73.800 77.200 ;
        RECT 76.600 76.800 77.000 77.200 ;
        RECT 73.400 75.200 73.700 76.800 ;
        RECT 69.400 74.800 69.800 75.200 ;
        RECT 72.600 74.800 73.000 75.200 ;
        RECT 73.400 74.800 73.800 75.200 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 75.800 75.100 76.200 75.200 ;
        RECT 75.000 74.800 76.200 75.100 ;
        RECT 76.600 74.800 77.000 75.200 ;
        RECT 67.800 73.800 68.200 74.200 ;
        RECT 67.800 73.200 68.100 73.800 ;
        RECT 67.800 72.800 68.200 73.200 ;
        RECT 69.400 69.200 69.700 74.800 ;
        RECT 70.200 73.800 70.600 74.200 ;
        RECT 70.200 73.200 70.500 73.800 ;
        RECT 70.200 72.800 70.600 73.200 ;
        RECT 72.600 69.800 73.000 70.200 ;
        RECT 76.600 70.100 76.900 74.800 ;
        RECT 77.400 71.200 77.700 85.800 ;
        RECT 78.200 81.800 78.600 82.200 ;
        RECT 78.200 79.200 78.500 81.800 ;
        RECT 79.000 79.200 79.300 85.800 ;
        RECT 80.600 84.800 81.000 85.200 ;
        RECT 80.600 84.200 80.900 84.800 ;
        RECT 80.600 83.800 81.000 84.200 ;
        RECT 81.400 82.100 81.700 96.800 ;
        RECT 82.200 92.100 82.600 97.900 ;
        RECT 87.800 97.800 88.200 98.200 ;
        RECT 83.000 93.800 83.400 94.200 ;
        RECT 83.000 93.200 83.300 93.800 ;
        RECT 83.000 92.800 83.400 93.200 ;
        RECT 83.800 93.100 84.200 95.900 ;
        RECT 85.400 91.800 85.800 92.200 ;
        RECT 88.600 92.100 89.000 97.900 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 91.800 94.800 92.200 95.200 ;
        RECT 83.000 88.800 83.400 89.200 ;
        RECT 83.800 89.100 84.200 89.200 ;
        RECT 84.600 89.100 85.000 89.200 ;
        RECT 83.800 88.800 85.000 89.100 ;
        RECT 83.000 87.200 83.300 88.800 ;
        RECT 85.400 88.200 85.700 91.800 ;
        RECT 91.000 89.200 91.300 94.800 ;
        RECT 91.000 88.800 91.400 89.200 ;
        RECT 85.400 87.800 85.800 88.200 ;
        RECT 80.600 81.800 81.700 82.100 ;
        RECT 82.200 86.800 82.600 87.200 ;
        RECT 83.000 86.800 83.400 87.200 ;
        RECT 84.600 86.800 85.000 87.200 ;
        RECT 78.200 78.800 78.600 79.200 ;
        RECT 79.000 78.800 79.400 79.200 ;
        RECT 80.600 75.200 80.900 81.800 ;
        RECT 82.200 75.200 82.500 86.800 ;
        RECT 83.000 86.200 83.300 86.800 ;
        RECT 83.000 85.800 83.400 86.200 ;
        RECT 84.600 85.200 84.900 86.800 ;
        RECT 91.800 86.200 92.100 94.800 ;
        RECT 92.600 94.200 92.900 101.800 ;
        RECT 94.200 98.800 94.600 99.200 ;
        RECT 92.600 93.800 93.000 94.200 ;
        RECT 91.800 85.800 92.200 86.200 ;
        RECT 84.600 84.800 85.000 85.200 ;
        RECT 83.000 77.800 83.400 78.200 ;
        RECT 80.600 74.800 81.000 75.200 ;
        RECT 82.200 74.800 82.600 75.200 ;
        RECT 78.200 73.800 78.600 74.200 ;
        RECT 78.200 72.200 78.500 73.800 ;
        RECT 78.200 71.800 78.600 72.200 ;
        RECT 77.400 70.800 77.800 71.200 ;
        RECT 76.600 69.800 77.700 70.100 ;
        RECT 67.000 68.800 67.400 69.200 ;
        RECT 69.400 68.800 69.800 69.200 ;
        RECT 67.000 68.200 67.300 68.800 ;
        RECT 67.000 67.800 67.400 68.200 ;
        RECT 67.800 66.800 68.200 67.200 ;
        RECT 68.600 67.100 69.000 67.200 ;
        RECT 68.600 66.800 69.700 67.100 ;
        RECT 67.800 66.200 68.100 66.800 ;
        RECT 59.800 65.800 60.200 66.200 ;
        RECT 62.200 65.800 62.600 66.200 ;
        RECT 66.200 65.800 66.600 66.200 ;
        RECT 67.800 65.800 68.200 66.200 ;
        RECT 59.800 65.200 60.100 65.800 ;
        RECT 59.800 64.800 60.200 65.200 ;
        RECT 60.600 63.800 61.000 64.200 ;
        RECT 58.200 55.800 58.600 56.200 ;
        RECT 58.200 47.200 58.500 55.800 ;
        RECT 59.000 52.100 59.400 57.900 ;
        RECT 59.800 48.800 60.200 49.200 ;
        RECT 59.800 48.200 60.100 48.800 ;
        RECT 59.800 47.800 60.200 48.200 ;
        RECT 60.600 47.200 60.900 63.800 ;
        RECT 62.200 56.200 62.500 65.800 ;
        RECT 66.200 59.100 66.600 59.200 ;
        RECT 67.000 59.100 67.400 59.200 ;
        RECT 66.200 58.800 67.400 59.100 ;
        RECT 62.200 55.800 62.600 56.200 ;
        RECT 62.200 54.800 62.600 55.200 ;
        RECT 61.400 53.800 61.800 54.200 ;
        RECT 61.400 53.200 61.700 53.800 ;
        RECT 61.400 52.800 61.800 53.200 ;
        RECT 61.400 48.200 61.700 52.800 ;
        RECT 62.200 52.200 62.500 54.800 ;
        RECT 62.200 51.800 62.600 52.200 ;
        RECT 63.800 52.100 64.200 57.900 ;
        RECT 65.400 53.100 65.800 55.900 ;
        RECT 66.200 54.800 66.600 55.200 ;
        RECT 64.600 51.800 65.000 52.200 ;
        RECT 64.600 49.200 64.900 51.800 ;
        RECT 64.600 48.800 65.000 49.200 ;
        RECT 61.400 47.800 61.800 48.200 ;
        RECT 58.200 46.800 58.600 47.200 ;
        RECT 60.600 46.800 61.000 47.200 ;
        RECT 64.600 47.100 65.000 47.200 ;
        RECT 65.400 47.100 65.800 47.200 ;
        RECT 64.600 46.800 65.800 47.100 ;
        RECT 66.200 46.200 66.500 54.800 ;
        RECT 67.800 54.100 68.200 54.200 ;
        RECT 68.600 54.100 69.000 54.200 ;
        RECT 67.800 53.800 69.000 54.100 ;
        RECT 69.400 53.200 69.700 66.800 ;
        RECT 70.200 65.100 70.600 67.900 ;
        RECT 71.800 63.100 72.200 68.900 ;
        RECT 72.600 68.200 72.900 69.800 ;
        RECT 72.600 67.800 73.000 68.200 ;
        RECT 73.400 66.100 73.800 66.200 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 73.400 65.800 74.600 66.100 ;
        RECT 76.600 63.100 77.000 68.900 ;
        RECT 71.800 61.800 72.200 62.200 ;
        RECT 71.800 59.200 72.100 61.800 ;
        RECT 77.400 60.200 77.700 69.800 ;
        RECT 79.000 69.100 79.400 69.200 ;
        RECT 79.800 69.100 80.200 69.200 ;
        RECT 79.000 68.800 80.200 69.100 ;
        RECT 77.400 59.800 77.800 60.200 ;
        RECT 71.800 58.800 72.200 59.200 ;
        RECT 73.400 55.800 73.800 56.200 ;
        RECT 73.400 55.200 73.700 55.800 ;
        RECT 70.200 54.800 70.600 55.200 ;
        RECT 73.400 54.800 73.800 55.200 ;
        RECT 74.200 54.800 74.600 55.200 ;
        RECT 78.200 54.800 78.600 55.200 ;
        RECT 79.000 54.800 79.400 55.200 ;
        RECT 70.200 54.200 70.500 54.800 ;
        RECT 70.200 53.800 70.600 54.200 ;
        RECT 67.000 53.100 67.400 53.200 ;
        RECT 67.800 53.100 68.200 53.200 ;
        RECT 67.000 52.800 68.200 53.100 ;
        RECT 68.600 52.800 69.000 53.200 ;
        RECT 69.400 52.800 69.800 53.200 ;
        RECT 72.600 53.100 73.000 53.200 ;
        RECT 73.400 53.100 73.800 53.200 ;
        RECT 72.600 52.800 73.800 53.100 ;
        RECT 68.600 49.200 68.900 52.800 ;
        RECT 68.600 48.800 69.000 49.200 ;
        RECT 68.600 46.800 69.000 47.200 ;
        RECT 68.600 46.200 68.900 46.800 ;
        RECT 57.400 45.800 57.800 46.200 ;
        RECT 58.200 45.800 58.600 46.200 ;
        RECT 59.800 45.800 60.200 46.200 ;
        RECT 63.000 46.100 63.400 46.200 ;
        RECT 63.800 46.100 64.200 46.200 ;
        RECT 63.000 45.800 64.200 46.100 ;
        RECT 66.200 45.800 66.600 46.200 ;
        RECT 68.600 45.800 69.000 46.200 ;
        RECT 57.400 44.200 57.700 45.800 ;
        RECT 57.400 43.800 57.800 44.200 ;
        RECT 58.200 43.100 58.500 45.800 ;
        RECT 57.400 42.800 58.500 43.100 ;
        RECT 57.400 35.200 57.700 42.800 ;
        RECT 59.800 39.200 60.100 45.800 ;
        RECT 59.800 38.800 60.200 39.200 ;
        RECT 65.400 38.800 65.800 39.200 ;
        RECT 65.400 38.200 65.700 38.800 ;
        RECT 65.400 37.800 65.800 38.200 ;
        RECT 64.600 36.800 65.000 37.200 ;
        RECT 64.600 36.200 64.900 36.800 ;
        RECT 64.600 35.800 65.000 36.200 ;
        RECT 65.400 36.100 65.800 36.200 ;
        RECT 66.200 36.100 66.600 36.200 ;
        RECT 65.400 35.800 66.600 36.100 ;
        RECT 67.800 35.800 68.200 36.200 ;
        RECT 57.400 34.800 57.800 35.200 ;
        RECT 58.200 35.100 58.600 35.200 ;
        RECT 59.000 35.100 59.400 35.200 ;
        RECT 58.200 34.800 59.400 35.100 ;
        RECT 57.400 29.200 57.700 34.800 ;
        RECT 67.800 33.200 68.100 35.800 ;
        RECT 69.400 35.200 69.700 52.800 ;
        RECT 71.000 45.100 71.400 47.900 ;
        RECT 71.800 47.800 72.200 48.200 ;
        RECT 71.800 47.200 72.100 47.800 ;
        RECT 71.800 46.800 72.200 47.200 ;
        RECT 71.800 44.800 72.200 45.200 ;
        RECT 71.800 39.200 72.100 44.800 ;
        RECT 72.600 43.100 73.000 48.900 ;
        RECT 71.800 38.800 72.200 39.200 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 71.800 35.100 72.200 35.200 ;
        RECT 72.600 35.100 73.000 35.200 ;
        RECT 71.800 34.800 73.000 35.100 ;
        RECT 69.400 34.200 69.700 34.800 ;
        RECT 69.400 33.800 69.800 34.200 ;
        RECT 59.000 33.100 59.400 33.200 ;
        RECT 59.800 33.100 60.200 33.200 ;
        RECT 59.000 32.800 60.200 33.100 ;
        RECT 67.800 32.800 68.200 33.200 ;
        RECT 68.600 32.800 69.000 33.200 ;
        RECT 63.800 31.800 64.200 32.200 ;
        RECT 57.400 28.800 57.800 29.200 ;
        RECT 63.800 28.200 64.100 31.800 ;
        RECT 65.400 29.800 65.800 30.200 ;
        RECT 65.400 29.200 65.700 29.800 ;
        RECT 68.600 29.200 68.900 32.800 ;
        RECT 69.400 32.200 69.700 33.800 ;
        RECT 69.400 31.800 69.800 32.200 ;
        RECT 64.600 28.800 65.000 29.200 ;
        RECT 65.400 28.800 65.800 29.200 ;
        RECT 67.800 28.800 68.200 29.200 ;
        RECT 68.600 28.800 69.000 29.200 ;
        RECT 63.800 27.800 64.200 28.200 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 62.200 27.100 62.600 27.200 ;
        RECT 61.400 26.800 62.600 27.100 ;
        RECT 63.800 25.800 64.200 26.200 ;
        RECT 59.800 24.100 60.200 24.200 ;
        RECT 60.600 24.100 61.000 24.200 ;
        RECT 59.800 23.800 61.000 24.100 ;
        RECT 61.400 22.800 61.800 23.200 ;
        RECT 60.600 15.800 61.000 16.200 ;
        RECT 60.600 15.200 60.900 15.800 ;
        RECT 57.400 15.100 57.800 15.200 ;
        RECT 56.600 14.800 57.800 15.100 ;
        RECT 60.600 14.800 61.000 15.200 ;
        RECT 57.400 14.200 57.700 14.800 ;
        RECT 55.800 13.800 56.200 14.200 ;
        RECT 57.400 13.800 57.800 14.200 ;
        RECT 59.000 14.100 59.400 14.200 ;
        RECT 59.800 14.100 60.200 14.200 ;
        RECT 59.000 13.800 60.200 14.100 ;
        RECT 55.800 13.200 56.100 13.800 ;
        RECT 61.400 13.200 61.700 22.800 ;
        RECT 63.000 13.800 63.400 14.200 ;
        RECT 55.800 12.800 56.200 13.200 ;
        RECT 59.000 13.100 59.400 13.200 ;
        RECT 59.800 13.100 60.200 13.200 ;
        RECT 61.400 13.100 61.800 13.200 ;
        RECT 59.000 12.800 60.200 13.100 ;
        RECT 60.600 12.800 61.800 13.100 ;
        RECT 60.600 9.200 60.900 12.800 ;
        RECT 47.000 6.100 47.400 6.200 ;
        RECT 47.800 6.100 48.200 6.200 ;
        RECT 47.000 5.800 48.200 6.100 ;
        RECT 50.200 5.800 50.600 6.200 ;
        RECT 51.000 5.800 51.400 6.200 ;
        RECT 51.800 5.100 52.200 7.900 ;
        RECT 52.600 7.800 53.000 8.200 ;
        RECT 52.600 7.200 52.900 7.800 ;
        RECT 52.600 6.800 53.000 7.200 ;
        RECT 53.400 3.100 53.800 8.900 ;
        RECT 55.000 6.100 55.400 6.200 ;
        RECT 55.800 6.100 56.200 6.200 ;
        RECT 55.000 5.800 56.200 6.100 ;
        RECT 58.200 3.100 58.600 8.900 ;
        RECT 60.600 8.800 61.000 9.200 ;
        RECT 63.000 6.200 63.300 13.800 ;
        RECT 63.800 9.200 64.100 25.800 ;
        RECT 64.600 25.200 64.900 28.800 ;
        RECT 67.800 28.200 68.100 28.800 ;
        RECT 67.800 27.800 68.200 28.200 ;
        RECT 74.200 26.200 74.500 54.800 ;
        RECT 75.800 52.800 76.200 53.200 ;
        RECT 75.000 51.800 75.400 52.200 ;
        RECT 75.000 46.200 75.300 51.800 ;
        RECT 75.000 45.800 75.400 46.200 ;
        RECT 75.800 35.200 76.100 52.800 ;
        RECT 76.600 47.800 77.000 48.200 ;
        RECT 76.600 47.200 76.900 47.800 ;
        RECT 76.600 46.800 77.000 47.200 ;
        RECT 77.400 43.100 77.800 48.900 ;
        RECT 78.200 42.200 78.500 54.800 ;
        RECT 79.000 52.200 79.300 54.800 ;
        RECT 79.800 53.800 80.200 54.200 ;
        RECT 79.000 51.800 79.400 52.200 ;
        RECT 79.800 49.200 80.100 53.800 ;
        RECT 80.600 52.200 80.900 74.800 ;
        RECT 83.000 74.200 83.300 77.800 ;
        RECT 84.600 75.200 84.900 84.800 ;
        RECT 87.000 83.800 87.400 84.200 ;
        RECT 83.800 74.800 84.200 75.200 ;
        RECT 84.600 74.800 85.000 75.200 ;
        RECT 81.400 73.800 81.800 74.200 ;
        RECT 82.200 73.800 82.600 74.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 81.400 72.200 81.700 73.800 ;
        RECT 81.400 71.800 81.800 72.200 ;
        RECT 81.400 66.800 81.800 67.200 ;
        RECT 81.400 66.200 81.700 66.800 ;
        RECT 81.400 65.800 81.800 66.200 ;
        RECT 82.200 59.200 82.500 73.800 ;
        RECT 82.200 58.800 82.600 59.200 ;
        RECT 83.000 58.100 83.300 73.800 ;
        RECT 83.800 61.200 84.100 74.800 ;
        RECT 85.400 72.100 85.800 72.200 ;
        RECT 86.200 72.100 86.600 72.200 ;
        RECT 85.400 71.800 86.600 72.100 ;
        RECT 84.600 70.800 85.000 71.200 ;
        RECT 84.600 66.200 84.900 70.800 ;
        RECT 87.000 69.200 87.300 83.800 ;
        RECT 91.000 78.800 91.400 79.200 ;
        RECT 88.600 72.100 89.000 77.900 ;
        RECT 91.000 75.200 91.300 78.800 ;
        RECT 91.800 76.200 92.100 85.800 ;
        RECT 91.800 75.800 92.200 76.200 ;
        RECT 91.000 74.800 91.400 75.200 ;
        RECT 92.600 74.200 92.900 93.800 ;
        RECT 93.400 92.100 93.800 97.900 ;
        RECT 93.400 88.100 93.800 88.200 ;
        RECT 94.200 88.100 94.500 98.800 ;
        RECT 95.800 96.200 96.100 113.800 ;
        RECT 96.600 113.200 96.900 114.800 ;
        RECT 98.200 114.200 98.500 125.800 ;
        RECT 99.000 123.200 99.300 125.800 ;
        RECT 99.800 125.100 100.200 125.200 ;
        RECT 100.600 125.100 101.000 125.200 ;
        RECT 99.800 124.800 101.000 125.100 ;
        RECT 102.200 124.200 102.500 125.800 ;
        RECT 103.800 124.800 104.200 125.200 ;
        RECT 102.200 123.800 102.600 124.200 ;
        RECT 99.000 122.800 99.400 123.200 ;
        RECT 99.000 117.100 99.400 117.200 ;
        RECT 99.800 117.100 100.200 117.200 ;
        RECT 99.000 116.800 100.200 117.100 ;
        RECT 98.200 113.800 98.600 114.200 ;
        RECT 99.000 113.800 99.400 114.200 ;
        RECT 96.600 112.800 97.000 113.200 ;
        RECT 97.400 111.800 97.800 112.200 ;
        RECT 97.400 108.200 97.700 111.800 ;
        RECT 99.000 111.200 99.300 113.800 ;
        RECT 101.400 111.800 101.800 112.200 ;
        RECT 102.200 112.100 102.600 117.900 ;
        RECT 99.000 110.800 99.400 111.200 ;
        RECT 99.000 109.800 99.400 110.200 ;
        RECT 97.400 107.800 97.800 108.200 ;
        RECT 99.000 106.200 99.300 109.800 ;
        RECT 101.400 107.200 101.700 111.800 ;
        RECT 103.800 109.200 104.100 124.800 ;
        RECT 110.200 123.100 110.600 128.900 ;
        RECT 113.400 126.200 113.700 131.800 ;
        RECT 115.000 131.200 115.300 134.800 ;
        RECT 115.800 134.200 116.100 134.800 ;
        RECT 115.800 133.800 116.200 134.200 ;
        RECT 116.600 133.100 117.000 135.900 ;
        RECT 118.200 132.100 118.600 137.900 ;
        RECT 119.000 134.200 119.300 146.800 ;
        RECT 123.800 143.100 124.200 148.900 ;
        RECT 124.600 146.800 125.000 147.200 ;
        RECT 124.600 146.200 124.900 146.800 ;
        RECT 124.600 145.800 125.000 146.200 ;
        RECT 127.000 145.800 127.400 146.200 ;
        RECT 127.000 145.200 127.300 145.800 ;
        RECT 127.000 144.800 127.400 145.200 ;
        RECT 120.600 142.100 121.000 142.200 ;
        RECT 121.400 142.100 121.800 142.200 ;
        RECT 120.600 141.800 121.800 142.100 ;
        RECT 127.800 139.200 128.100 154.800 ;
        RECT 128.600 154.200 128.900 154.800 ;
        RECT 128.600 153.800 129.000 154.200 ;
        RECT 129.400 151.200 129.700 154.800 ;
        RECT 133.400 154.200 133.700 154.800 ;
        RECT 133.400 153.800 133.800 154.200 ;
        RECT 135.000 152.800 135.400 153.200 ;
        RECT 135.000 152.200 135.300 152.800 ;
        RECT 135.000 151.800 135.400 152.200 ;
        RECT 129.400 150.800 129.800 151.200 ;
        RECT 135.800 151.100 136.100 164.800 ;
        RECT 139.800 162.100 140.200 168.900 ;
        RECT 140.600 162.100 141.000 168.900 ;
        RECT 141.400 163.100 141.800 168.900 ;
        RECT 142.200 166.800 142.600 167.200 ;
        RECT 142.200 166.200 142.500 166.800 ;
        RECT 142.200 165.800 142.600 166.200 ;
        RECT 143.000 163.100 143.400 168.900 ;
        RECT 143.800 168.800 144.200 169.200 ;
        RECT 143.800 168.200 144.100 168.800 ;
        RECT 143.800 167.800 144.200 168.200 ;
        RECT 144.600 163.100 145.000 168.900 ;
        RECT 145.400 162.100 145.800 168.900 ;
        RECT 146.200 162.100 146.600 168.900 ;
        RECT 147.000 162.100 147.400 168.900 ;
        RECT 150.200 166.800 150.600 167.200 ;
        RECT 137.400 153.100 137.800 155.900 ;
        RECT 139.000 152.100 139.400 157.900 ;
        RECT 139.800 155.800 140.200 156.200 ;
        RECT 139.800 155.100 140.100 155.800 ;
        RECT 139.800 154.700 140.200 155.100 ;
        RECT 139.800 152.800 140.200 153.200 ;
        RECT 142.200 152.800 142.600 153.200 ;
        RECT 135.000 150.800 136.100 151.100 ;
        RECT 128.600 143.100 129.000 148.900 ;
        RECT 130.200 145.100 130.600 147.900 ;
        RECT 131.000 147.800 131.400 148.200 ;
        RECT 131.000 147.200 131.300 147.800 ;
        RECT 131.000 146.800 131.400 147.200 ;
        RECT 134.200 146.800 134.600 147.200 ;
        RECT 134.200 146.200 134.500 146.800 ;
        RECT 135.000 146.200 135.300 150.800 ;
        RECT 139.800 148.200 140.100 152.800 ;
        RECT 139.800 147.800 140.200 148.200 ;
        RECT 131.000 146.100 131.400 146.200 ;
        RECT 131.800 146.100 132.200 146.200 ;
        RECT 131.000 145.800 132.200 146.100 ;
        RECT 132.600 145.800 133.000 146.200 ;
        RECT 134.200 145.800 134.600 146.200 ;
        RECT 135.000 145.800 135.400 146.200 ;
        RECT 135.800 146.100 136.200 146.200 ;
        RECT 136.600 146.100 137.000 146.200 ;
        RECT 135.800 145.800 137.000 146.100 ;
        RECT 127.800 138.800 128.200 139.200 ;
        RECT 119.800 134.800 120.200 135.200 ;
        RECT 119.800 134.200 120.100 134.800 ;
        RECT 119.000 133.800 119.400 134.200 ;
        RECT 119.800 133.800 120.200 134.200 ;
        RECT 119.000 133.200 119.300 133.800 ;
        RECT 119.000 132.800 119.400 133.200 ;
        RECT 123.000 132.100 123.400 137.900 ;
        RECT 127.800 135.200 128.100 138.800 ;
        RECT 131.800 136.100 132.100 145.800 ;
        RECT 132.600 145.200 132.900 145.800 ;
        RECT 132.600 144.800 133.000 145.200 ;
        RECT 132.600 136.800 133.000 137.200 ;
        RECT 132.600 136.100 132.900 136.800 ;
        RECT 131.800 135.800 132.900 136.100 ;
        RECT 132.600 135.200 132.900 135.800 ;
        RECT 134.200 135.800 134.600 136.200 ;
        RECT 134.200 135.200 134.500 135.800 ;
        RECT 126.200 135.100 126.600 135.200 ;
        RECT 127.000 135.100 127.400 135.200 ;
        RECT 126.200 134.800 127.400 135.100 ;
        RECT 127.800 134.800 128.200 135.200 ;
        RECT 130.200 135.100 130.600 135.200 ;
        RECT 131.000 135.100 131.400 135.200 ;
        RECT 130.200 134.800 131.400 135.100 ;
        RECT 131.800 134.800 132.200 135.200 ;
        RECT 132.600 134.800 133.000 135.200 ;
        RECT 134.200 134.800 134.600 135.200 ;
        RECT 127.800 134.100 128.200 134.200 ;
        RECT 128.600 134.100 129.000 134.200 ;
        RECT 127.800 133.800 129.000 134.100 ;
        RECT 123.800 132.800 124.200 133.200 ;
        RECT 115.000 130.800 115.400 131.200 ;
        RECT 116.600 129.100 117.000 129.200 ;
        RECT 117.400 129.100 117.800 129.200 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 114.200 123.800 114.600 124.200 ;
        RECT 104.600 115.100 105.000 115.200 ;
        RECT 105.400 115.100 105.800 115.200 ;
        RECT 104.600 114.800 105.800 115.100 ;
        RECT 105.400 113.800 105.800 114.200 ;
        RECT 103.800 108.800 104.200 109.200 ;
        RECT 99.800 106.800 100.200 107.200 ;
        RECT 101.400 106.800 101.800 107.200 ;
        RECT 103.000 106.800 103.400 107.200 ;
        RECT 99.800 106.200 100.100 106.800 ;
        RECT 103.000 106.200 103.300 106.800 ;
        RECT 99.000 105.800 99.400 106.200 ;
        RECT 99.800 105.800 100.200 106.200 ;
        RECT 100.600 105.800 101.000 106.200 ;
        RECT 102.200 105.800 102.600 106.200 ;
        RECT 103.000 105.800 103.400 106.200 ;
        RECT 104.600 105.800 105.000 106.200 ;
        RECT 100.600 104.200 100.900 105.800 ;
        RECT 100.600 103.800 101.000 104.200 ;
        RECT 96.600 101.800 97.000 102.200 ;
        RECT 96.600 99.200 96.900 101.800 ;
        RECT 96.600 98.800 97.000 99.200 ;
        RECT 99.800 99.100 100.200 99.200 ;
        RECT 100.600 99.100 101.000 99.200 ;
        RECT 99.800 98.800 101.000 99.100 ;
        RECT 99.800 96.800 100.200 97.200 ;
        RECT 99.800 96.200 100.100 96.800 ;
        RECT 95.000 93.100 95.400 95.900 ;
        RECT 95.800 95.800 96.200 96.200 ;
        RECT 96.600 96.100 97.000 96.200 ;
        RECT 97.400 96.100 97.800 96.200 ;
        RECT 96.600 95.800 97.800 96.100 ;
        RECT 99.800 95.800 100.200 96.200 ;
        RECT 95.800 93.800 96.200 94.200 ;
        RECT 96.600 93.800 97.000 94.200 ;
        RECT 98.200 93.800 98.600 94.200 ;
        RECT 95.800 93.200 96.100 93.800 ;
        RECT 93.400 87.800 94.500 88.100 ;
        RECT 95.800 92.800 96.200 93.200 ;
        RECT 95.000 86.800 95.400 87.200 ;
        RECT 95.000 86.200 95.300 86.800 ;
        RECT 95.800 86.200 96.100 92.800 ;
        RECT 96.600 89.200 96.900 93.800 ;
        RECT 98.200 93.200 98.500 93.800 ;
        RECT 98.200 92.800 98.600 93.200 ;
        RECT 99.800 91.800 100.200 92.200 ;
        RECT 99.800 90.200 100.100 91.800 ;
        RECT 99.800 89.800 100.200 90.200 ;
        RECT 96.600 88.800 97.000 89.200 ;
        RECT 102.200 88.200 102.500 105.800 ;
        RECT 103.800 101.800 104.200 102.200 ;
        RECT 103.000 92.100 103.400 97.900 ;
        RECT 103.800 89.100 104.100 101.800 ;
        RECT 104.600 97.200 104.900 105.800 ;
        RECT 104.600 96.800 105.000 97.200 ;
        RECT 104.600 94.800 105.000 95.200 ;
        RECT 104.600 94.200 104.900 94.800 ;
        RECT 105.400 94.200 105.700 113.800 ;
        RECT 107.000 112.100 107.400 117.900 ;
        RECT 112.600 116.800 113.000 117.200 ;
        RECT 112.600 116.200 112.900 116.800 ;
        RECT 107.800 113.800 108.200 114.200 ;
        RECT 107.800 113.200 108.100 113.800 ;
        RECT 107.800 112.800 108.200 113.200 ;
        RECT 108.600 113.100 109.000 115.900 ;
        RECT 112.600 115.800 113.000 116.200 ;
        RECT 114.200 115.200 114.500 123.800 ;
        RECT 115.000 123.100 115.400 128.900 ;
        RECT 116.600 128.800 117.800 129.100 ;
        RECT 115.800 127.800 116.200 128.200 ;
        RECT 115.800 127.200 116.100 127.800 ;
        RECT 115.800 126.800 116.200 127.200 ;
        RECT 116.600 125.100 117.000 127.900 ;
        RECT 119.800 123.100 120.200 128.900 ;
        RECT 123.800 128.200 124.100 132.800 ;
        RECT 129.400 130.800 129.800 131.200 ;
        RECT 120.600 127.800 121.000 128.200 ;
        RECT 123.800 127.800 124.200 128.200 ;
        RECT 120.600 127.200 120.900 127.800 ;
        RECT 120.600 126.800 121.000 127.200 ;
        RECT 123.800 126.800 124.200 127.200 ;
        RECT 123.800 126.300 124.100 126.800 ;
        RECT 123.800 125.900 124.200 126.300 ;
        RECT 124.600 123.100 125.000 128.900 ;
        RECT 127.000 128.800 127.400 129.200 ;
        RECT 127.000 128.200 127.300 128.800 ;
        RECT 126.200 125.100 126.600 127.900 ;
        RECT 127.000 127.800 127.400 128.200 ;
        RECT 127.000 127.100 127.400 127.200 ;
        RECT 127.800 127.100 128.200 127.200 ;
        RECT 127.000 126.800 128.200 127.100 ;
        RECT 129.400 126.200 129.700 130.800 ;
        RECT 131.000 130.200 131.300 134.800 ;
        RECT 131.800 133.200 132.100 134.800 ;
        RECT 135.000 133.200 135.300 145.800 ;
        RECT 141.400 143.100 141.800 148.900 ;
        RECT 135.800 135.100 136.200 135.200 ;
        RECT 135.800 134.800 136.900 135.100 ;
        RECT 131.800 132.800 132.200 133.200 ;
        RECT 135.000 132.800 135.400 133.200 ;
        RECT 131.000 129.800 131.400 130.200 ;
        RECT 130.200 128.100 130.600 128.200 ;
        RECT 131.000 128.100 131.400 128.200 ;
        RECT 130.200 127.800 131.400 128.100 ;
        RECT 136.600 127.200 136.900 134.800 ;
        RECT 137.400 134.800 137.800 135.200 ;
        RECT 131.800 126.800 132.200 127.200 ;
        RECT 133.400 126.800 133.800 127.200 ;
        RECT 134.200 126.800 134.600 127.200 ;
        RECT 135.000 127.100 135.400 127.200 ;
        RECT 135.800 127.100 136.200 127.200 ;
        RECT 135.000 126.800 136.200 127.100 ;
        RECT 136.600 126.800 137.000 127.200 ;
        RECT 131.800 126.200 132.100 126.800 ;
        RECT 128.600 125.800 129.000 126.200 ;
        RECT 129.400 125.800 129.800 126.200 ;
        RECT 131.800 125.800 132.200 126.200 ;
        RECT 128.600 123.200 128.900 125.800 ;
        RECT 129.400 123.200 129.700 125.800 ;
        RECT 133.400 124.200 133.700 126.800 ;
        RECT 134.200 126.200 134.500 126.800 ;
        RECT 137.400 126.200 137.700 134.800 ;
        RECT 139.000 131.800 139.400 132.200 ;
        RECT 140.600 131.800 141.000 132.200 ;
        RECT 141.400 132.100 141.800 137.900 ;
        RECT 139.000 128.200 139.300 131.800 ;
        RECT 139.000 127.800 139.400 128.200 ;
        RECT 140.600 127.200 140.900 131.800 ;
        RECT 142.200 129.200 142.500 152.800 ;
        RECT 143.800 152.100 144.200 157.900 ;
        RECT 145.400 152.100 145.800 152.200 ;
        RECT 146.200 152.100 146.600 152.200 ;
        RECT 145.400 151.800 146.600 152.100 ;
        RECT 150.200 149.200 150.500 166.800 ;
        RECT 155.800 165.100 156.200 167.900 ;
        RECT 156.600 167.800 157.000 168.200 ;
        RECT 156.600 167.200 156.900 167.800 ;
        RECT 156.600 166.800 157.000 167.200 ;
        RECT 151.800 161.800 152.200 162.200 ;
        RECT 144.600 145.800 145.000 146.200 ;
        RECT 144.600 145.200 144.900 145.800 ;
        RECT 144.600 144.800 145.000 145.200 ;
        RECT 146.200 143.100 146.600 148.900 ;
        RECT 150.200 148.800 150.600 149.200 ;
        RECT 151.800 148.200 152.100 161.800 ;
        RECT 155.800 158.800 156.200 159.200 ;
        RECT 154.200 152.800 154.600 153.200 ;
        RECT 152.600 151.800 153.000 152.200 ;
        RECT 147.000 147.800 147.400 148.200 ;
        RECT 147.000 147.200 147.300 147.800 ;
        RECT 147.000 146.800 147.400 147.200 ;
        RECT 143.800 135.100 144.200 135.200 ;
        RECT 144.600 135.100 145.000 135.200 ;
        RECT 143.800 134.800 145.000 135.100 ;
        RECT 143.000 132.800 143.400 133.200 ;
        RECT 142.200 128.800 142.600 129.200 ;
        RECT 143.000 128.200 143.300 132.800 ;
        RECT 146.200 132.100 146.600 137.900 ;
        RECT 147.000 134.200 147.300 146.800 ;
        RECT 147.800 145.100 148.200 147.900 ;
        RECT 151.800 147.800 152.200 148.200 ;
        RECT 152.600 147.200 152.900 151.800 ;
        RECT 154.200 147.200 154.500 152.800 ;
        RECT 155.000 151.800 155.400 152.200 ;
        RECT 155.000 148.200 155.300 151.800 ;
        RECT 155.800 150.200 156.100 158.800 ;
        RECT 156.600 152.200 156.900 166.800 ;
        RECT 157.400 163.100 157.800 168.900 ;
        RECT 159.000 166.100 159.400 166.200 ;
        RECT 159.800 166.100 160.200 166.200 ;
        RECT 159.000 165.800 160.200 166.100 ;
        RECT 162.200 163.100 162.600 168.900 ;
        RECT 165.400 165.800 165.800 166.200 ;
        RECT 166.200 166.100 166.600 166.200 ;
        RECT 167.000 166.100 167.400 166.200 ;
        RECT 166.200 165.800 167.400 166.100 ;
        RECT 168.600 165.800 169.000 166.200 ;
        RECT 170.200 165.800 170.600 166.200 ;
        RECT 171.000 165.800 171.400 166.200 ;
        RECT 172.600 166.100 173.000 166.200 ;
        RECT 173.400 166.100 173.800 166.200 ;
        RECT 172.600 165.800 173.800 166.100 ;
        RECT 174.200 165.800 174.600 166.200 ;
        RECT 176.600 166.100 177.000 166.200 ;
        RECT 177.400 166.100 177.800 166.200 ;
        RECT 176.600 165.800 177.800 166.100 ;
        RECT 164.600 161.800 165.000 162.200 ;
        RECT 164.600 161.200 164.900 161.800 ;
        RECT 165.400 161.200 165.700 165.800 ;
        RECT 168.600 164.200 168.900 165.800 ;
        RECT 170.200 165.200 170.500 165.800 ;
        RECT 170.200 164.800 170.600 165.200 ;
        RECT 168.600 163.800 169.000 164.200 ;
        RECT 167.800 161.800 168.200 162.200 ;
        RECT 164.600 160.800 165.000 161.200 ;
        RECT 165.400 160.800 165.800 161.200 ;
        RECT 158.200 153.800 158.600 154.200 ;
        RECT 156.600 151.800 157.000 152.200 ;
        RECT 155.800 149.800 156.200 150.200 ;
        RECT 155.800 148.200 156.100 149.800 ;
        RECT 158.200 149.200 158.500 153.800 ;
        RECT 159.800 152.100 160.200 158.900 ;
        RECT 160.600 152.100 161.000 158.900 ;
        RECT 161.400 152.100 161.800 157.900 ;
        RECT 162.200 153.800 162.600 154.200 ;
        RECT 162.200 153.200 162.500 153.800 ;
        RECT 162.200 152.800 162.600 153.200 ;
        RECT 163.000 152.100 163.400 157.900 ;
        RECT 163.800 152.800 164.200 153.200 ;
        RECT 163.800 152.200 164.100 152.800 ;
        RECT 163.800 151.800 164.200 152.200 ;
        RECT 164.600 152.100 165.000 157.900 ;
        RECT 165.400 152.100 165.800 158.900 ;
        RECT 166.200 152.100 166.600 158.900 ;
        RECT 167.000 152.100 167.400 158.900 ;
        RECT 167.800 152.200 168.100 161.800 ;
        RECT 171.000 156.200 171.300 165.800 ;
        RECT 172.600 161.800 173.000 162.200 ;
        RECT 172.600 156.200 172.900 161.800 ;
        RECT 171.000 155.800 171.400 156.200 ;
        RECT 172.600 155.800 173.000 156.200 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 167.800 151.800 168.200 152.200 ;
        RECT 171.800 151.800 172.200 152.200 ;
        RECT 161.400 150.800 161.800 151.200 ;
        RECT 158.200 148.800 158.600 149.200 ;
        RECT 161.400 148.200 161.700 150.800 ;
        RECT 163.800 148.200 164.100 151.800 ;
        RECT 171.800 151.200 172.100 151.800 ;
        RECT 171.800 150.800 172.200 151.200 ;
        RECT 173.400 150.200 173.700 154.800 ;
        RECT 173.400 149.800 173.800 150.200 ;
        RECT 155.000 147.800 155.400 148.200 ;
        RECT 155.800 147.800 156.200 148.200 ;
        RECT 161.400 147.800 161.800 148.200 ;
        RECT 163.800 147.800 164.200 148.200 ;
        RECT 149.400 146.800 149.800 147.200 ;
        RECT 152.600 146.800 153.000 147.200 ;
        RECT 154.200 146.800 154.600 147.200 ;
        RECT 156.600 147.100 157.000 147.200 ;
        RECT 157.400 147.100 157.800 147.200 ;
        RECT 156.600 146.800 157.800 147.100 ;
        RECT 148.600 145.800 149.000 146.200 ;
        RECT 148.600 145.200 148.900 145.800 ;
        RECT 148.600 144.800 149.000 145.200 ;
        RECT 149.400 143.200 149.700 146.800 ;
        RECT 154.200 146.100 154.600 146.200 ;
        RECT 155.000 146.100 155.400 146.200 ;
        RECT 154.200 145.800 155.400 146.100 ;
        RECT 156.600 145.800 157.000 146.200 ;
        RECT 159.800 145.800 160.200 146.200 ;
        RECT 156.600 145.200 156.900 145.800 ;
        RECT 156.600 144.800 157.000 145.200 ;
        RECT 149.400 142.800 149.800 143.200 ;
        RECT 154.200 141.800 154.600 142.200 ;
        RECT 148.600 137.800 149.000 138.200 ;
        RECT 148.600 136.200 148.900 137.800 ;
        RECT 147.000 133.800 147.400 134.200 ;
        RECT 147.800 133.100 148.200 135.900 ;
        RECT 148.600 135.800 149.000 136.200 ;
        RECT 151.000 133.800 151.400 134.200 ;
        RECT 153.400 133.800 153.800 134.200 ;
        RECT 148.600 131.800 149.000 132.200 ;
        RECT 147.800 130.800 148.200 131.200 ;
        RECT 147.800 129.200 148.100 130.800 ;
        RECT 147.800 128.800 148.200 129.200 ;
        RECT 143.000 127.800 143.400 128.200 ;
        RECT 148.600 127.200 148.900 131.800 ;
        RECT 151.000 131.200 151.300 133.800 ;
        RECT 151.800 132.800 152.200 133.200 ;
        RECT 151.000 130.800 151.400 131.200 ;
        RECT 151.800 129.200 152.100 132.800 ;
        RECT 150.200 129.100 150.600 129.200 ;
        RECT 151.000 129.100 151.400 129.200 ;
        RECT 150.200 128.800 151.400 129.100 ;
        RECT 151.800 128.800 152.200 129.200 ;
        RECT 149.400 128.100 149.800 128.200 ;
        RECT 150.200 128.100 150.600 128.200 ;
        RECT 149.400 127.800 150.600 128.100 ;
        RECT 140.600 126.800 141.000 127.200 ;
        RECT 147.000 126.800 147.400 127.200 ;
        RECT 148.600 126.800 149.000 127.200 ;
        RECT 147.000 126.200 147.300 126.800 ;
        RECT 134.200 125.800 134.600 126.200 ;
        RECT 135.800 125.800 136.200 126.200 ;
        RECT 137.400 125.800 137.800 126.200 ;
        RECT 140.600 125.800 141.000 126.200 ;
        RECT 147.000 125.800 147.400 126.200 ;
        RECT 135.800 125.200 136.100 125.800 ;
        RECT 135.800 124.800 136.200 125.200 ;
        RECT 133.400 123.800 133.800 124.200 ;
        RECT 128.600 122.800 129.000 123.200 ;
        RECT 129.400 122.800 129.800 123.200 ;
        RECT 133.400 122.800 133.800 123.200 ;
        RECT 114.200 114.800 114.600 115.200 ;
        RECT 115.000 114.800 115.400 115.200 ;
        RECT 109.400 112.800 109.800 113.200 ;
        RECT 109.400 112.200 109.700 112.800 ;
        RECT 109.400 111.800 109.800 112.200 ;
        RECT 107.000 110.800 107.400 111.200 ;
        RECT 107.000 109.200 107.300 110.800 ;
        RECT 107.000 108.800 107.400 109.200 ;
        RECT 109.400 108.800 109.800 109.200 ;
        RECT 110.200 109.100 110.600 109.200 ;
        RECT 111.000 109.100 111.400 109.200 ;
        RECT 110.200 108.800 111.400 109.100 ;
        RECT 109.400 108.200 109.700 108.800 ;
        RECT 109.400 107.800 109.800 108.200 ;
        RECT 106.200 106.800 106.600 107.200 ;
        RECT 107.000 107.100 107.400 107.200 ;
        RECT 107.800 107.100 108.200 107.200 ;
        RECT 107.000 106.800 108.200 107.100 ;
        RECT 106.200 95.200 106.500 106.800 ;
        RECT 109.400 106.200 109.700 107.800 ;
        RECT 109.400 105.800 109.800 106.200 ;
        RECT 112.600 105.800 113.000 106.200 ;
        RECT 110.200 101.800 110.600 102.200 ;
        RECT 106.200 94.800 106.600 95.200 ;
        RECT 104.600 93.800 105.000 94.200 ;
        RECT 105.400 93.800 105.800 94.200 ;
        RECT 106.200 93.800 106.600 94.200 ;
        RECT 103.800 88.800 104.900 89.100 ;
        RECT 101.400 87.800 101.800 88.200 ;
        RECT 102.200 87.800 102.600 88.200 ;
        RECT 101.400 87.200 101.700 87.800 ;
        RECT 99.000 86.800 99.400 87.200 ;
        RECT 101.400 86.800 101.800 87.200 ;
        RECT 99.000 86.200 99.300 86.800 ;
        RECT 93.400 85.800 93.800 86.200 ;
        RECT 95.000 85.800 95.400 86.200 ;
        RECT 95.800 85.800 96.200 86.200 ;
        RECT 97.400 86.100 97.800 86.200 ;
        RECT 98.200 86.100 98.600 86.200 ;
        RECT 97.400 85.800 98.600 86.100 ;
        RECT 99.000 85.800 99.400 86.200 ;
        RECT 99.800 85.800 100.200 86.200 ;
        RECT 102.200 85.800 102.600 86.200 ;
        RECT 103.000 85.800 103.400 86.200 ;
        RECT 93.400 84.200 93.700 85.800 ;
        RECT 95.000 85.200 95.300 85.800 ;
        RECT 95.000 84.800 95.400 85.200 ;
        RECT 93.400 83.800 93.800 84.200 ;
        RECT 92.600 73.800 93.000 74.200 ;
        RECT 92.600 69.200 92.900 73.800 ;
        RECT 93.400 72.100 93.800 77.900 ;
        RECT 95.000 73.100 95.400 75.900 ;
        RECT 95.800 74.200 96.100 85.800 ;
        RECT 96.600 83.800 97.000 84.200 ;
        RECT 96.600 79.200 96.900 83.800 ;
        RECT 96.600 78.800 97.000 79.200 ;
        RECT 97.400 77.800 97.800 78.200 ;
        RECT 97.400 76.200 97.700 77.800 ;
        RECT 97.400 75.800 97.800 76.200 ;
        RECT 99.800 75.200 100.100 85.800 ;
        RECT 100.600 81.800 101.000 82.200 ;
        RECT 100.600 80.200 100.900 81.800 ;
        RECT 100.600 79.800 101.000 80.200 ;
        RECT 100.600 79.200 100.900 79.800 ;
        RECT 102.200 79.200 102.500 85.800 ;
        RECT 103.000 80.100 103.300 85.800 ;
        RECT 103.800 85.100 104.200 87.900 ;
        RECT 103.000 79.800 104.100 80.100 ;
        RECT 100.600 78.800 101.000 79.200 ;
        RECT 102.200 78.800 102.600 79.200 ;
        RECT 100.600 76.800 101.000 77.200 ;
        RECT 100.600 75.200 100.900 76.800 ;
        RECT 99.800 74.800 100.200 75.200 ;
        RECT 100.600 74.800 101.000 75.200 ;
        RECT 95.800 74.100 96.200 74.200 ;
        RECT 96.600 74.100 97.000 74.200 ;
        RECT 95.800 73.800 97.000 74.100 ;
        RECT 97.400 74.100 97.800 74.200 ;
        RECT 98.200 74.100 98.600 74.200 ;
        RECT 97.400 73.800 98.600 74.100 ;
        RECT 97.400 71.800 97.800 72.200 ;
        RECT 95.000 70.800 95.400 71.200 ;
        RECT 87.000 68.800 87.400 69.200 ;
        RECT 91.000 68.800 91.400 69.200 ;
        RECT 92.600 68.800 93.000 69.200 ;
        RECT 91.000 68.200 91.300 68.800 ;
        RECT 91.000 67.800 91.400 68.200 ;
        RECT 91.000 67.200 91.300 67.800 ;
        RECT 85.400 67.100 85.800 67.200 ;
        RECT 86.200 67.100 86.600 67.200 ;
        RECT 85.400 66.800 86.600 67.100 ;
        RECT 91.000 66.800 91.400 67.200 ;
        RECT 84.600 65.800 85.000 66.200 ;
        RECT 85.400 65.800 85.800 66.200 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 89.400 65.800 89.800 66.200 ;
        RECT 84.600 64.200 84.900 65.800 ;
        RECT 85.400 65.200 85.700 65.800 ;
        RECT 86.200 65.200 86.500 65.800 ;
        RECT 85.400 64.800 85.800 65.200 ;
        RECT 86.200 64.800 86.600 65.200 ;
        RECT 84.600 63.800 85.000 64.200 ;
        RECT 85.400 61.200 85.700 64.800 ;
        RECT 89.400 62.200 89.700 65.800 ;
        RECT 91.800 64.800 92.200 65.200 ;
        RECT 89.400 61.800 89.800 62.200 ;
        RECT 83.800 60.800 84.200 61.200 ;
        RECT 85.400 60.800 85.800 61.200 ;
        RECT 83.800 59.800 84.200 60.200 ;
        RECT 83.800 59.200 84.100 59.800 ;
        RECT 83.800 58.800 84.200 59.200 ;
        RECT 82.200 57.800 83.300 58.100 ;
        RECT 82.200 54.200 82.500 57.800 ;
        RECT 83.000 54.800 83.400 55.200 ;
        RECT 81.400 54.100 81.800 54.200 ;
        RECT 82.200 54.100 82.600 54.200 ;
        RECT 81.400 53.800 82.600 54.100 ;
        RECT 80.600 51.800 81.000 52.200 ;
        RECT 79.800 48.800 80.200 49.200 ;
        RECT 80.600 45.100 81.000 47.900 ;
        RECT 81.400 46.800 81.800 47.200 ;
        RECT 81.400 46.200 81.700 46.800 ;
        RECT 81.400 45.800 81.800 46.200 ;
        RECT 81.400 44.800 81.800 45.200 ;
        RECT 81.400 43.200 81.700 44.800 ;
        RECT 81.400 42.800 81.800 43.200 ;
        RECT 82.200 43.100 82.600 48.900 ;
        RECT 78.200 41.800 78.600 42.200 ;
        RECT 75.800 34.800 76.200 35.200 ;
        RECT 77.400 34.800 77.800 35.200 ;
        RECT 75.800 33.200 76.100 34.800 ;
        RECT 77.400 34.200 77.700 34.800 ;
        RECT 77.400 33.800 77.800 34.200 ;
        RECT 75.800 32.800 76.200 33.200 ;
        RECT 77.400 32.800 77.800 33.200 ;
        RECT 75.800 31.800 76.200 32.200 ;
        RECT 75.800 29.200 76.100 31.800 ;
        RECT 75.800 28.800 76.200 29.200 ;
        RECT 76.600 27.800 77.000 28.200 ;
        RECT 76.600 27.200 76.900 27.800 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 77.400 26.200 77.700 32.800 ;
        RECT 74.200 25.800 74.600 26.200 ;
        RECT 75.000 25.800 75.400 26.200 ;
        RECT 77.400 25.800 77.800 26.200 ;
        RECT 64.600 24.800 65.000 25.200 ;
        RECT 67.800 24.800 68.200 25.200 ;
        RECT 67.000 16.800 67.400 17.200 ;
        RECT 67.000 15.200 67.300 16.800 ;
        RECT 67.800 16.200 68.100 24.800 ;
        RECT 75.000 24.200 75.300 25.800 ;
        RECT 75.000 23.800 75.400 24.200 ;
        RECT 68.600 21.800 69.000 22.200 ;
        RECT 68.600 19.200 68.900 21.800 ;
        RECT 75.000 19.800 75.400 20.200 ;
        RECT 68.600 18.800 69.000 19.200 ;
        RECT 67.800 16.100 68.200 16.200 ;
        RECT 68.600 16.100 69.000 16.200 ;
        RECT 67.800 15.800 69.000 16.100 ;
        RECT 75.000 15.200 75.300 19.800 ;
        RECT 78.200 19.200 78.500 41.800 ;
        RECT 81.400 39.200 81.700 42.800 ;
        RECT 80.600 38.800 81.000 39.200 ;
        RECT 81.400 38.800 81.800 39.200 ;
        RECT 79.000 38.100 79.400 38.200 ;
        RECT 79.800 38.100 80.200 38.200 ;
        RECT 79.000 37.800 80.200 38.100 ;
        RECT 80.600 35.200 80.900 38.800 ;
        RECT 83.000 36.200 83.300 54.800 ;
        RECT 86.200 52.100 86.600 57.900 ;
        RECT 90.200 54.700 90.600 55.100 ;
        RECT 88.600 54.100 89.000 54.200 ;
        RECT 87.800 53.800 89.000 54.100 ;
        RECT 87.800 52.200 88.100 53.800 ;
        RECT 90.200 53.200 90.500 54.700 ;
        RECT 90.200 52.800 90.600 53.200 ;
        RECT 87.800 51.800 88.200 52.200 ;
        RECT 91.000 52.100 91.400 57.900 ;
        RECT 91.800 56.200 92.100 64.800 ;
        RECT 94.200 63.100 94.600 68.900 ;
        RECT 91.800 55.800 92.200 56.200 ;
        RECT 83.800 46.800 84.200 47.200 ;
        RECT 83.800 46.200 84.100 46.800 ;
        RECT 83.800 45.800 84.200 46.200 ;
        RECT 87.000 43.100 87.400 48.900 ;
        RECT 87.800 44.200 88.100 51.800 ;
        RECT 90.200 49.100 90.600 49.200 ;
        RECT 91.000 49.100 91.400 49.200 ;
        RECT 90.200 48.800 91.400 49.100 ;
        RECT 91.800 46.200 92.100 55.800 ;
        RECT 92.600 53.100 93.000 55.900 ;
        RECT 95.000 55.200 95.300 70.800 ;
        RECT 97.400 55.200 97.700 71.800 ;
        RECT 99.800 71.200 100.100 74.800 ;
        RECT 100.600 73.800 101.000 74.200 ;
        RECT 100.600 73.200 100.900 73.800 ;
        RECT 100.600 72.800 101.000 73.200 ;
        RECT 102.200 73.100 102.600 73.200 ;
        RECT 103.000 73.100 103.400 73.200 ;
        RECT 102.200 72.800 103.400 73.100 ;
        RECT 101.400 71.800 101.800 72.200 ;
        RECT 99.800 70.800 100.200 71.200 ;
        RECT 101.400 69.200 101.700 71.800 ;
        RECT 103.800 71.200 104.100 79.800 ;
        RECT 104.600 75.200 104.900 88.800 ;
        RECT 105.400 83.100 105.800 88.900 ;
        RECT 106.200 88.200 106.500 93.800 ;
        RECT 107.800 92.100 108.200 97.900 ;
        RECT 109.400 93.100 109.800 95.900 ;
        RECT 110.200 95.200 110.500 101.800 ;
        RECT 112.600 99.200 112.900 105.800 ;
        RECT 113.400 103.100 113.800 108.900 ;
        RECT 114.200 99.200 114.500 114.800 ;
        RECT 115.000 114.200 115.300 114.800 ;
        RECT 115.000 113.800 115.400 114.200 ;
        RECT 115.000 112.100 115.400 112.200 ;
        RECT 115.800 112.100 116.200 112.200 ;
        RECT 118.200 112.100 118.600 117.900 ;
        RECT 121.400 115.800 121.800 116.200 ;
        RECT 121.400 115.200 121.700 115.800 ;
        RECT 121.400 114.800 121.800 115.200 ;
        RECT 121.400 113.800 121.800 114.200 ;
        RECT 121.400 113.200 121.700 113.800 ;
        RECT 121.400 112.800 121.800 113.200 ;
        RECT 115.000 111.800 116.200 112.100 ;
        RECT 115.800 106.100 116.200 106.200 ;
        RECT 116.600 106.100 117.000 106.200 ;
        RECT 115.800 105.800 117.000 106.100 ;
        RECT 118.200 103.100 118.600 108.900 ;
        RECT 119.800 105.100 120.200 107.900 ;
        RECT 120.600 105.100 121.000 107.900 ;
        RECT 121.400 107.200 121.700 112.800 ;
        RECT 123.000 112.100 123.400 117.900 ;
        RECT 124.600 113.100 125.000 115.900 ;
        RECT 132.600 115.800 133.000 116.200 ;
        RECT 132.600 115.200 132.900 115.800 ;
        RECT 133.400 115.200 133.700 122.800 ;
        RECT 132.600 114.800 133.000 115.200 ;
        RECT 133.400 114.800 133.800 115.200 ;
        RECT 126.200 111.800 126.600 112.200 ;
        RECT 121.400 106.800 121.800 107.200 ;
        RECT 120.600 103.800 121.000 104.200 ;
        RECT 112.600 98.800 113.000 99.200 ;
        RECT 114.200 98.800 114.600 99.200 ;
        RECT 110.200 94.800 110.600 95.200 ;
        RECT 112.600 95.100 113.000 95.200 ;
        RECT 113.400 95.100 113.800 95.200 ;
        RECT 112.600 94.800 113.800 95.100 ;
        RECT 114.200 94.800 114.600 95.200 ;
        RECT 115.000 94.800 115.400 95.200 ;
        RECT 106.200 87.800 106.600 88.200 ;
        RECT 106.200 86.800 106.600 87.200 ;
        RECT 106.200 86.300 106.500 86.800 ;
        RECT 106.200 85.900 106.600 86.300 ;
        RECT 110.200 83.100 110.600 88.900 ;
        RECT 114.200 84.200 114.500 94.800 ;
        RECT 115.000 94.200 115.300 94.800 ;
        RECT 115.000 93.800 115.400 94.200 ;
        RECT 115.000 92.800 115.400 93.200 ;
        RECT 117.400 93.100 117.800 93.200 ;
        RECT 118.200 93.100 118.600 93.200 ;
        RECT 117.400 92.800 118.600 93.100 ;
        RECT 115.000 88.200 115.300 92.800 ;
        RECT 115.800 91.800 116.200 92.200 ;
        RECT 115.800 89.200 116.100 91.800 ;
        RECT 120.600 89.200 120.900 103.800 ;
        RECT 122.200 103.100 122.600 108.900 ;
        RECT 126.200 107.200 126.500 111.800 ;
        RECT 126.200 106.800 126.600 107.200 ;
        RECT 123.000 105.900 123.400 106.300 ;
        RECT 126.200 106.200 126.500 106.800 ;
        RECT 123.000 104.200 123.300 105.900 ;
        RECT 126.200 105.800 126.600 106.200 ;
        RECT 123.000 103.800 123.400 104.200 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 115.800 88.800 116.200 89.200 ;
        RECT 120.600 88.800 121.000 89.200 ;
        RECT 115.000 87.800 115.400 88.200 ;
        RECT 116.600 86.800 117.000 87.200 ;
        RECT 116.600 86.200 116.900 86.800 ;
        RECT 122.200 86.200 122.500 94.800 ;
        RECT 123.000 92.100 123.400 98.900 ;
        RECT 123.800 92.100 124.200 98.900 ;
        RECT 124.600 92.100 125.000 98.900 ;
        RECT 125.400 92.100 125.800 97.900 ;
        RECT 126.200 93.200 126.500 105.800 ;
        RECT 127.000 103.100 127.400 108.900 ;
        RECT 130.200 105.100 130.600 107.900 ;
        RECT 131.000 106.800 131.400 107.200 ;
        RECT 131.000 106.200 131.300 106.800 ;
        RECT 131.000 105.800 131.400 106.200 ;
        RECT 131.800 103.100 132.200 108.900 ;
        RECT 128.600 102.100 129.000 102.200 ;
        RECT 129.400 102.100 129.800 102.200 ;
        RECT 128.600 101.800 129.800 102.100 ;
        RECT 133.400 101.200 133.700 114.800 ;
        RECT 135.800 114.100 136.200 114.200 ;
        RECT 136.600 114.100 137.000 114.200 ;
        RECT 135.800 113.800 137.000 114.100 ;
        RECT 135.800 112.800 136.200 113.200 ;
        RECT 134.200 107.800 134.600 108.200 ;
        RECT 134.200 106.200 134.500 107.800 ;
        RECT 135.800 107.200 136.100 112.800 ;
        RECT 137.400 112.200 137.700 125.800 ;
        RECT 140.600 122.200 140.900 125.800 ;
        RECT 152.600 123.100 153.000 128.900 ;
        RECT 153.400 126.200 153.700 133.800 ;
        RECT 154.200 133.200 154.500 141.800 ;
        RECT 159.800 138.200 160.100 145.800 ;
        RECT 163.000 144.800 163.400 145.200 ;
        RECT 163.000 139.200 163.300 144.800 ;
        RECT 166.200 142.100 166.600 148.900 ;
        RECT 167.000 142.100 167.400 148.900 ;
        RECT 167.800 143.100 168.200 148.900 ;
        RECT 168.600 146.800 169.000 147.200 ;
        RECT 168.600 146.200 168.900 146.800 ;
        RECT 168.600 145.800 169.000 146.200 ;
        RECT 169.400 143.100 169.800 148.900 ;
        RECT 170.200 148.800 170.600 149.200 ;
        RECT 170.200 148.200 170.500 148.800 ;
        RECT 170.200 147.800 170.600 148.200 ;
        RECT 171.000 143.100 171.400 148.900 ;
        RECT 170.200 141.800 170.600 142.200 ;
        RECT 171.800 142.100 172.200 148.900 ;
        RECT 172.600 142.100 173.000 148.900 ;
        RECT 173.400 142.100 173.800 148.900 ;
        RECT 174.200 142.200 174.500 165.800 ;
        RECT 177.400 154.800 177.800 155.200 ;
        RECT 176.600 152.800 177.000 153.200 ;
        RECT 175.800 151.800 176.200 152.200 ;
        RECT 175.000 147.800 175.400 148.200 ;
        RECT 174.200 141.800 174.600 142.200 ;
        RECT 163.000 138.800 163.400 139.200 ;
        RECT 159.800 137.800 160.200 138.200 ;
        RECT 163.800 137.800 164.200 138.200 ;
        RECT 156.600 136.800 157.000 137.200 ;
        RECT 156.600 135.200 156.900 136.800 ;
        RECT 163.800 136.200 164.100 137.800 ;
        RECT 168.600 136.800 169.000 137.200 ;
        RECT 159.800 135.800 160.200 136.200 ;
        RECT 163.000 135.800 163.400 136.200 ;
        RECT 163.800 135.800 164.200 136.200 ;
        RECT 166.200 135.800 166.600 136.200 ;
        RECT 156.600 134.800 157.000 135.200 ;
        RECT 157.400 134.800 157.800 135.200 ;
        RECT 157.400 134.200 157.700 134.800 ;
        RECT 159.800 134.200 160.100 135.800 ;
        RECT 163.000 135.200 163.300 135.800 ;
        RECT 160.600 135.100 161.000 135.200 ;
        RECT 160.600 134.800 161.700 135.100 ;
        RECT 163.000 134.800 163.400 135.200 ;
        RECT 157.400 133.800 157.800 134.200 ;
        RECT 159.800 133.800 160.200 134.200 ;
        RECT 154.200 132.800 154.600 133.200 ;
        RECT 159.800 132.800 160.200 133.200 ;
        RECT 159.800 132.200 160.100 132.800 ;
        RECT 155.000 131.800 155.400 132.200 ;
        RECT 159.800 131.800 160.200 132.200 ;
        RECT 155.000 126.200 155.300 131.800 ;
        RECT 160.600 129.800 161.000 130.200 ;
        RECT 155.800 126.800 156.200 127.200 ;
        RECT 153.400 125.800 153.800 126.200 ;
        RECT 155.000 125.800 155.400 126.200 ;
        RECT 140.600 121.800 141.000 122.200 ;
        RECT 139.000 117.100 139.400 117.200 ;
        RECT 139.800 117.100 140.200 117.200 ;
        RECT 139.000 116.800 140.200 117.100 ;
        RECT 137.400 111.800 137.800 112.200 ;
        RECT 143.000 112.100 143.400 117.900 ;
        RECT 143.800 114.800 144.200 115.200 ;
        RECT 146.200 114.800 146.600 115.200 ;
        RECT 143.800 113.200 144.100 114.800 ;
        RECT 146.200 114.200 146.500 114.800 ;
        RECT 146.200 113.800 146.600 114.200 ;
        RECT 143.800 112.800 144.200 113.200 ;
        RECT 144.600 112.800 145.000 113.200 ;
        RECT 135.800 106.800 136.200 107.200 ;
        RECT 134.200 105.800 134.600 106.200 ;
        RECT 135.000 102.800 135.400 103.200 ;
        RECT 136.600 103.100 137.000 108.900 ;
        RECT 143.800 107.800 144.200 108.200 ;
        RECT 143.800 107.200 144.100 107.800 ;
        RECT 143.000 106.800 143.400 107.200 ;
        RECT 143.800 106.800 144.200 107.200 ;
        RECT 143.000 106.200 143.300 106.800 ;
        RECT 143.000 105.800 143.400 106.200 ;
        RECT 143.800 105.800 144.200 106.200 ;
        RECT 143.800 105.200 144.100 105.800 ;
        RECT 143.800 104.800 144.200 105.200 ;
        RECT 133.400 100.800 133.800 101.200 ;
        RECT 133.400 99.200 133.700 100.800 ;
        RECT 126.200 92.800 126.600 93.200 ;
        RECT 123.800 90.800 124.200 91.200 ;
        RECT 123.800 88.200 124.100 90.800 ;
        RECT 126.200 90.100 126.500 92.800 ;
        RECT 127.000 92.100 127.400 97.900 ;
        RECT 127.800 93.800 128.200 94.200 ;
        RECT 127.800 92.200 128.100 93.800 ;
        RECT 127.800 91.800 128.200 92.200 ;
        RECT 128.600 92.100 129.000 97.900 ;
        RECT 129.400 92.100 129.800 98.900 ;
        RECT 130.200 92.100 130.600 98.900 ;
        RECT 133.400 98.800 133.800 99.200 ;
        RECT 126.200 89.800 127.300 90.100 ;
        RECT 123.800 87.800 124.200 88.200 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 117.400 85.800 117.800 86.200 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 121.400 86.100 121.800 86.200 ;
        RECT 120.600 85.800 121.800 86.100 ;
        RECT 122.200 86.100 122.600 86.200 ;
        RECT 123.000 86.100 123.400 86.200 ;
        RECT 122.200 85.800 123.400 86.100 ;
        RECT 117.400 85.200 117.700 85.800 ;
        RECT 119.000 85.200 119.300 85.800 ;
        RECT 115.800 84.800 116.200 85.200 ;
        RECT 117.400 84.800 117.800 85.200 ;
        RECT 119.000 84.800 119.400 85.200 ;
        RECT 114.200 83.800 114.600 84.200 ;
        RECT 114.200 81.800 114.600 82.200 ;
        RECT 114.200 79.200 114.500 81.800 ;
        RECT 115.800 79.200 116.100 84.800 ;
        RECT 120.600 81.200 120.900 85.800 ;
        RECT 123.000 85.100 123.400 85.200 ;
        RECT 123.800 85.100 124.200 85.200 ;
        RECT 124.600 85.100 125.000 87.900 ;
        RECT 125.400 85.800 125.800 86.200 ;
        RECT 123.000 84.800 124.200 85.100 ;
        RECT 120.600 80.800 121.000 81.200 ;
        RECT 111.000 78.800 111.400 79.200 ;
        RECT 114.200 78.800 114.600 79.200 ;
        RECT 115.800 78.800 116.200 79.200 ;
        RECT 105.400 77.800 105.800 78.200 ;
        RECT 108.600 77.800 109.000 78.200 ;
        RECT 105.400 75.200 105.700 77.800 ;
        RECT 108.600 75.200 108.900 77.800 ;
        RECT 111.000 75.200 111.300 78.800 ;
        RECT 113.400 78.100 113.800 78.200 ;
        RECT 114.200 78.100 114.600 78.200 ;
        RECT 113.400 77.800 114.600 78.100 ;
        RECT 113.400 77.100 113.800 77.200 ;
        RECT 112.600 76.800 113.800 77.100 ;
        RECT 118.200 76.800 118.600 77.200 ;
        RECT 112.600 76.200 112.900 76.800 ;
        RECT 112.600 75.800 113.000 76.200 ;
        RECT 118.200 75.200 118.500 76.800 ;
        RECT 104.600 74.800 105.000 75.200 ;
        RECT 105.400 74.800 105.800 75.200 ;
        RECT 106.200 75.100 106.600 75.200 ;
        RECT 107.000 75.100 107.400 75.200 ;
        RECT 106.200 74.800 107.400 75.100 ;
        RECT 108.600 74.800 109.000 75.200 ;
        RECT 111.000 74.800 111.400 75.200 ;
        RECT 118.200 74.800 118.600 75.200 ;
        RECT 104.600 72.800 105.000 73.200 ;
        RECT 103.800 70.800 104.200 71.200 ;
        RECT 98.200 68.800 98.600 69.200 ;
        RECT 98.200 68.200 98.500 68.800 ;
        RECT 98.200 67.800 98.600 68.200 ;
        RECT 98.200 66.800 98.600 67.200 ;
        RECT 98.200 66.300 98.500 66.800 ;
        RECT 98.200 65.900 98.600 66.300 ;
        RECT 99.000 63.100 99.400 68.900 ;
        RECT 99.800 68.800 100.200 69.200 ;
        RECT 101.400 68.800 101.800 69.200 ;
        RECT 98.200 59.800 98.600 60.200 ;
        RECT 94.200 55.100 94.600 55.200 ;
        RECT 95.000 55.100 95.400 55.200 ;
        RECT 94.200 54.800 95.400 55.100 ;
        RECT 97.400 54.800 97.800 55.200 ;
        RECT 95.800 54.100 96.200 54.200 ;
        RECT 96.600 54.100 97.000 54.200 ;
        RECT 95.800 53.800 97.000 54.100 ;
        RECT 98.200 53.200 98.500 59.800 ;
        RECT 99.800 55.200 100.100 68.800 ;
        RECT 100.600 65.100 101.000 67.900 ;
        RECT 101.400 67.800 101.800 68.200 ;
        RECT 101.400 67.200 101.700 67.800 ;
        RECT 101.400 66.800 101.800 67.200 ;
        RECT 103.000 67.100 103.400 67.200 ;
        RECT 103.800 67.100 104.200 67.200 ;
        RECT 103.000 66.800 104.200 67.100 ;
        RECT 103.800 62.800 104.200 63.200 ;
        RECT 100.600 59.800 101.000 60.200 ;
        RECT 100.600 59.200 100.900 59.800 ;
        RECT 100.600 58.800 101.000 59.200 ;
        RECT 100.600 57.800 101.000 58.200 ;
        RECT 99.000 54.800 99.400 55.200 ;
        RECT 99.800 54.800 100.200 55.200 ;
        RECT 96.600 53.100 97.000 53.200 ;
        RECT 97.400 53.100 97.800 53.200 ;
        RECT 96.600 52.800 97.800 53.100 ;
        RECT 98.200 52.800 98.600 53.200 ;
        RECT 97.400 48.800 97.800 49.200 ;
        RECT 97.400 48.200 97.700 48.800 ;
        RECT 92.600 47.800 93.000 48.200 ;
        RECT 93.400 47.800 93.800 48.200 ;
        RECT 97.400 48.100 97.800 48.200 ;
        RECT 98.200 48.100 98.600 48.200 ;
        RECT 97.400 47.800 98.600 48.100 ;
        RECT 99.000 48.100 99.300 54.800 ;
        RECT 99.800 54.200 100.100 54.800 ;
        RECT 99.800 53.800 100.200 54.200 ;
        RECT 100.600 49.200 100.900 57.800 ;
        RECT 103.000 52.100 103.400 57.900 ;
        RECT 103.000 50.800 103.400 51.200 ;
        RECT 100.600 48.800 101.000 49.200 ;
        RECT 99.000 47.800 100.100 48.100 ;
        RECT 92.600 46.200 92.900 47.800 ;
        RECT 93.400 47.200 93.700 47.800 ;
        RECT 93.400 46.800 93.800 47.200 ;
        RECT 99.000 46.800 99.400 47.200 ;
        RECT 91.800 45.800 92.200 46.200 ;
        RECT 92.600 45.800 93.000 46.200 ;
        RECT 97.400 46.100 97.800 46.200 ;
        RECT 98.200 46.100 98.600 46.200 ;
        RECT 97.400 45.800 98.600 46.100 ;
        RECT 87.800 43.800 88.200 44.200 ;
        RECT 89.400 43.800 89.800 44.200 ;
        RECT 83.800 36.800 84.200 37.200 ;
        RECT 83.800 36.200 84.100 36.800 ;
        RECT 83.000 35.800 83.400 36.200 ;
        RECT 83.800 35.800 84.200 36.200 ;
        RECT 79.800 34.800 80.200 35.200 ;
        RECT 80.600 34.800 81.000 35.200 ;
        RECT 82.200 35.100 82.600 35.200 ;
        RECT 83.000 35.100 83.400 35.200 ;
        RECT 82.200 34.800 83.400 35.100 ;
        RECT 87.000 34.800 87.400 35.200 ;
        RECT 79.800 33.200 80.100 34.800 ;
        RECT 83.800 33.800 84.200 34.200 ;
        RECT 85.400 33.800 85.800 34.200 ;
        RECT 79.800 32.800 80.200 33.200 ;
        RECT 81.400 33.100 81.800 33.200 ;
        RECT 82.200 33.100 82.600 33.200 ;
        RECT 81.400 32.800 82.600 33.100 ;
        RECT 79.000 31.800 79.400 32.200 ;
        RECT 78.200 18.800 78.600 19.200 ;
        RECT 79.000 16.200 79.300 31.800 ;
        RECT 79.800 29.200 80.100 32.800 ;
        RECT 79.800 28.800 80.200 29.200 ;
        RECT 82.200 29.100 82.600 29.200 ;
        RECT 83.000 29.100 83.400 29.200 ;
        RECT 82.200 28.800 83.400 29.100 ;
        RECT 79.800 26.800 80.200 27.200 ;
        RECT 79.800 26.200 80.100 26.800 ;
        RECT 79.800 25.800 80.200 26.200 ;
        RECT 79.800 19.100 80.200 19.200 ;
        RECT 80.600 19.100 81.000 19.200 ;
        RECT 79.800 18.800 81.000 19.100 ;
        RECT 79.000 15.800 79.400 16.200 ;
        RECT 65.400 15.100 65.800 15.200 ;
        RECT 66.200 15.100 66.600 15.200 ;
        RECT 65.400 14.800 66.600 15.100 ;
        RECT 67.000 14.800 67.400 15.200 ;
        RECT 71.800 14.800 72.200 15.200 ;
        RECT 75.000 14.800 75.400 15.200 ;
        RECT 71.800 14.200 72.100 14.800 ;
        RECT 69.400 13.800 69.800 14.200 ;
        RECT 71.800 13.800 72.200 14.200 ;
        RECT 73.400 14.100 73.800 14.200 ;
        RECT 74.200 14.100 74.600 14.200 ;
        RECT 73.400 13.800 74.600 14.100 ;
        RECT 69.400 9.200 69.700 13.800 ;
        RECT 73.400 11.800 73.800 12.200 ;
        RECT 82.200 12.100 82.600 17.900 ;
        RECT 83.000 13.800 83.400 14.200 ;
        RECT 63.800 8.800 64.200 9.200 ;
        RECT 65.400 9.100 65.800 9.200 ;
        RECT 66.200 9.100 66.600 9.200 ;
        RECT 65.400 8.800 66.600 9.100 ;
        RECT 63.000 5.800 63.400 6.200 ;
        RECT 67.800 3.100 68.200 8.900 ;
        RECT 69.400 8.800 69.800 9.200 ;
        RECT 71.800 6.800 72.200 7.200 ;
        RECT 71.800 6.300 72.100 6.800 ;
        RECT 71.800 5.900 72.200 6.300 ;
        RECT 72.600 3.100 73.000 8.900 ;
        RECT 73.400 6.200 73.700 11.800 ;
        RECT 73.400 5.800 73.800 6.200 ;
        RECT 74.200 5.100 74.600 7.900 ;
        RECT 75.000 5.100 75.400 7.900 ;
        RECT 76.600 3.100 77.000 8.900 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 78.200 7.200 78.500 7.800 ;
        RECT 78.200 6.800 78.600 7.200 ;
        RECT 77.400 6.100 77.800 6.200 ;
        RECT 78.200 6.100 78.600 6.200 ;
        RECT 77.400 5.800 78.600 6.100 ;
        RECT 81.400 3.100 81.800 8.900 ;
        RECT 83.000 7.200 83.300 13.800 ;
        RECT 83.800 9.200 84.100 33.800 ;
        RECT 85.400 32.200 85.700 33.800 ;
        RECT 87.000 33.200 87.300 34.800 ;
        RECT 87.800 34.200 88.100 43.800 ;
        RECT 88.600 36.800 89.000 37.200 ;
        RECT 88.600 35.200 88.900 36.800 ;
        RECT 89.400 35.200 89.700 43.800 ;
        RECT 91.800 37.200 92.100 45.800 ;
        RECT 91.800 36.800 92.200 37.200 ;
        RECT 91.000 35.800 91.400 36.200 ;
        RECT 91.000 35.200 91.300 35.800 ;
        RECT 88.600 34.800 89.000 35.200 ;
        RECT 89.400 34.800 89.800 35.200 ;
        RECT 91.000 34.800 91.400 35.200 ;
        RECT 87.800 33.800 88.200 34.200 ;
        RECT 87.000 32.800 87.400 33.200 ;
        RECT 85.400 31.800 85.800 32.200 ;
        RECT 84.600 23.100 85.000 28.900 ;
        RECT 87.800 27.200 88.100 33.800 ;
        RECT 92.600 29.200 92.900 45.800 ;
        RECT 99.000 39.200 99.300 46.800 ;
        RECT 94.200 38.800 94.600 39.200 ;
        RECT 99.000 38.800 99.400 39.200 ;
        RECT 94.200 33.200 94.500 38.800 ;
        RECT 94.200 32.800 94.600 33.200 ;
        RECT 95.000 33.100 95.400 35.900 ;
        RECT 95.800 34.800 96.200 35.200 ;
        RECT 95.800 34.200 96.100 34.800 ;
        RECT 95.800 33.800 96.200 34.200 ;
        RECT 96.600 32.100 97.000 37.900 ;
        RECT 97.400 35.800 97.800 36.200 ;
        RECT 97.400 35.100 97.700 35.800 ;
        RECT 97.400 34.700 97.800 35.100 ;
        RECT 87.800 26.800 88.200 27.200 ;
        RECT 88.600 26.800 89.000 27.200 ;
        RECT 86.200 15.800 86.600 16.200 ;
        RECT 86.200 15.100 86.500 15.800 ;
        RECT 86.200 14.700 86.600 15.100 ;
        RECT 87.000 12.100 87.400 17.900 ;
        RECT 87.800 17.200 88.100 26.800 ;
        RECT 88.600 26.300 88.900 26.800 ;
        RECT 88.600 25.900 89.000 26.300 ;
        RECT 89.400 23.100 89.800 28.900 ;
        RECT 91.800 28.800 92.200 29.200 ;
        RECT 92.600 28.800 93.000 29.200 ;
        RECT 91.800 28.200 92.100 28.800 ;
        RECT 91.000 25.100 91.400 27.900 ;
        RECT 91.800 27.800 92.200 28.200 ;
        RECT 95.000 27.100 95.400 27.200 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 95.000 26.800 96.200 27.100 ;
        RECT 99.800 26.200 100.100 47.800 ;
        RECT 101.400 47.800 101.800 48.200 ;
        RECT 101.400 47.200 101.700 47.800 ;
        RECT 100.600 46.800 101.000 47.200 ;
        RECT 101.400 46.800 101.800 47.200 ;
        RECT 100.600 43.200 100.900 46.800 ;
        RECT 103.000 46.200 103.300 50.800 ;
        RECT 103.800 49.200 104.100 62.800 ;
        RECT 103.800 48.800 104.200 49.200 ;
        RECT 104.600 48.200 104.900 72.800 ;
        RECT 105.400 65.200 105.700 74.800 ;
        RECT 106.200 73.800 106.600 74.200 ;
        RECT 110.200 73.800 110.600 74.200 ;
        RECT 112.600 74.100 113.000 74.200 ;
        RECT 114.200 74.100 114.600 74.200 ;
        RECT 112.600 73.800 114.600 74.100 ;
        RECT 115.800 74.100 116.200 74.200 ;
        RECT 118.200 74.100 118.600 74.200 ;
        RECT 115.800 73.800 118.600 74.100 ;
        RECT 106.200 66.200 106.500 73.800 ;
        RECT 110.200 72.200 110.500 73.800 ;
        RECT 115.800 72.800 116.200 73.200 ;
        RECT 119.000 72.800 119.400 73.200 ;
        RECT 107.800 71.800 108.200 72.200 ;
        RECT 110.200 71.800 110.600 72.200 ;
        RECT 107.800 69.200 108.100 71.800 ;
        RECT 110.200 69.800 110.600 70.200 ;
        RECT 107.800 68.800 108.200 69.200 ;
        RECT 107.000 66.800 107.400 67.200 ;
        RECT 107.000 66.200 107.300 66.800 ;
        RECT 106.200 65.800 106.600 66.200 ;
        RECT 107.000 65.800 107.400 66.200 ;
        RECT 105.400 64.800 105.800 65.200 ;
        RECT 106.200 64.200 106.500 65.800 ;
        RECT 107.800 65.100 108.200 67.900 ;
        RECT 106.200 63.800 106.600 64.200 ;
        RECT 109.400 63.100 109.800 68.900 ;
        RECT 110.200 68.200 110.500 69.800 ;
        RECT 111.000 68.800 111.400 69.200 ;
        RECT 115.800 69.100 116.100 72.800 ;
        RECT 119.000 72.200 119.300 72.800 ;
        RECT 119.000 71.800 119.400 72.200 ;
        RECT 118.200 70.800 118.600 71.200 ;
        RECT 118.200 69.200 118.500 70.800 ;
        RECT 116.600 69.100 117.000 69.200 ;
        RECT 110.200 67.800 110.600 68.200 ;
        RECT 111.000 66.200 111.300 68.800 ;
        RECT 111.000 65.800 111.400 66.200 ;
        RECT 114.200 63.100 114.600 68.900 ;
        RECT 115.800 68.800 117.000 69.100 ;
        RECT 118.200 68.800 118.600 69.200 ;
        RECT 116.600 68.100 117.000 68.200 ;
        RECT 117.400 68.100 117.800 68.200 ;
        RECT 116.600 67.800 117.800 68.100 ;
        RECT 117.400 66.800 117.800 67.200 ;
        RECT 115.800 64.800 116.200 65.200 ;
        RECT 110.200 59.800 110.600 60.200 ;
        RECT 106.200 55.000 106.600 55.100 ;
        RECT 107.000 55.000 107.400 55.100 ;
        RECT 106.200 54.700 107.400 55.000 ;
        RECT 105.400 53.800 105.800 54.200 ;
        RECT 105.400 52.200 105.700 53.800 ;
        RECT 105.400 51.800 105.800 52.200 ;
        RECT 107.800 52.100 108.200 57.900 ;
        RECT 109.400 53.100 109.800 55.900 ;
        RECT 110.200 53.200 110.500 59.800 ;
        RECT 115.000 56.800 115.400 57.200 ;
        RECT 115.000 55.200 115.300 56.800 ;
        RECT 115.800 55.200 116.100 64.800 ;
        RECT 117.400 59.200 117.700 66.800 ;
        RECT 120.600 66.200 120.900 80.800 ;
        RECT 123.800 78.200 124.100 84.800 ;
        RECT 122.200 77.800 122.600 78.200 ;
        RECT 123.800 77.800 124.200 78.200 ;
        RECT 122.200 75.200 122.500 77.800 ;
        RECT 123.000 77.100 123.400 77.200 ;
        RECT 123.800 77.100 124.200 77.200 ;
        RECT 123.000 76.800 124.200 77.100 ;
        RECT 124.600 76.800 125.000 77.200 ;
        RECT 122.200 74.800 122.600 75.200 ;
        RECT 123.800 74.800 124.200 75.200 ;
        RECT 121.400 73.800 121.800 74.200 ;
        RECT 121.400 68.200 121.700 73.800 ;
        RECT 123.800 71.200 124.100 74.800 ;
        RECT 124.600 74.200 124.900 76.800 ;
        RECT 125.400 75.200 125.700 85.800 ;
        RECT 126.200 83.100 126.600 88.900 ;
        RECT 127.000 88.200 127.300 89.800 ;
        RECT 127.000 87.800 127.400 88.200 ;
        RECT 127.800 85.800 128.200 86.200 ;
        RECT 127.800 81.200 128.100 85.800 ;
        RECT 131.000 83.100 131.400 88.900 ;
        RECT 135.000 87.200 135.300 102.800 ;
        RECT 137.400 93.800 137.800 94.200 ;
        RECT 135.800 91.800 136.200 92.200 ;
        RECT 135.800 89.200 136.100 91.800 ;
        RECT 135.800 88.800 136.200 89.200 ;
        RECT 135.000 86.800 135.400 87.200 ;
        RECT 137.400 86.200 137.700 93.800 ;
        RECT 140.600 92.100 141.000 98.900 ;
        RECT 141.400 92.100 141.800 98.900 ;
        RECT 142.200 92.100 142.600 97.900 ;
        RECT 143.000 93.800 143.400 94.200 ;
        RECT 143.000 92.200 143.300 93.800 ;
        RECT 143.000 91.800 143.400 92.200 ;
        RECT 143.800 92.100 144.200 97.900 ;
        RECT 144.600 93.200 144.900 112.800 ;
        RECT 147.000 111.800 147.400 112.200 ;
        RECT 147.800 112.100 148.200 117.900 ;
        RECT 149.400 113.100 149.800 115.900 ;
        RECT 151.000 112.800 151.400 113.200 ;
        RECT 151.800 113.100 152.200 115.900 ;
        RECT 152.600 113.800 153.000 114.200 ;
        RECT 152.600 113.200 152.900 113.800 ;
        RECT 152.600 112.800 153.000 113.200 ;
        RECT 151.000 112.200 151.300 112.800 ;
        RECT 150.200 111.800 150.600 112.200 ;
        RECT 151.000 111.800 151.400 112.200 ;
        RECT 153.400 112.100 153.800 117.900 ;
        RECT 155.000 114.800 155.400 115.200 ;
        RECT 155.000 113.200 155.300 114.800 ;
        RECT 155.000 112.800 155.400 113.200 ;
        RECT 146.200 106.800 146.600 107.200 ;
        RECT 146.200 106.200 146.500 106.800 ;
        RECT 147.000 106.200 147.300 111.800 ;
        RECT 147.800 107.800 148.200 108.200 ;
        RECT 147.800 107.200 148.100 107.800 ;
        RECT 147.800 106.800 148.200 107.200 ;
        RECT 149.400 106.800 149.800 107.200 ;
        RECT 146.200 105.800 146.600 106.200 ;
        RECT 147.000 105.800 147.400 106.200 ;
        RECT 147.800 106.100 148.200 106.200 ;
        RECT 148.600 106.100 149.000 106.200 ;
        RECT 147.800 105.800 149.000 106.100 ;
        RECT 147.000 101.200 147.300 105.800 ;
        RECT 149.400 104.200 149.700 106.800 ;
        RECT 149.400 103.800 149.800 104.200 ;
        RECT 147.000 100.800 147.400 101.200 ;
        RECT 144.600 92.800 145.000 93.200 ;
        RECT 140.600 90.800 141.000 91.200 ;
        RECT 140.600 88.200 140.900 90.800 ;
        RECT 144.600 88.200 144.900 92.800 ;
        RECT 145.400 92.100 145.800 97.900 ;
        RECT 146.200 92.100 146.600 98.900 ;
        RECT 147.000 92.100 147.400 98.900 ;
        RECT 147.800 92.100 148.200 98.900 ;
        RECT 150.200 90.100 150.500 111.800 ;
        RECT 151.800 103.100 152.200 108.900 ;
        RECT 155.800 108.200 156.100 126.800 ;
        RECT 157.400 123.100 157.800 128.900 ;
        RECT 159.000 125.100 159.400 127.900 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 159.800 124.200 160.100 126.800 ;
        RECT 160.600 126.200 160.900 129.800 ;
        RECT 161.400 127.200 161.700 134.800 ;
        RECT 163.000 127.800 163.400 128.200 ;
        RECT 163.000 127.200 163.300 127.800 ;
        RECT 163.800 127.200 164.100 135.800 ;
        RECT 166.200 135.200 166.500 135.800 ;
        RECT 168.600 135.200 168.900 136.800 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 167.000 135.100 167.400 135.200 ;
        RECT 167.800 135.100 168.200 135.200 ;
        RECT 167.000 134.800 168.200 135.100 ;
        RECT 168.600 134.800 169.000 135.200 ;
        RECT 167.000 133.800 167.400 134.200 ;
        RECT 167.000 133.200 167.300 133.800 ;
        RECT 167.000 132.800 167.400 133.200 ;
        RECT 167.800 132.800 168.200 133.200 ;
        RECT 164.600 127.800 165.000 128.200 ;
        RECT 167.000 127.800 167.400 128.200 ;
        RECT 161.400 126.800 161.800 127.200 ;
        RECT 163.000 126.800 163.400 127.200 ;
        RECT 163.800 126.800 164.200 127.200 ;
        RECT 164.600 126.200 164.900 127.800 ;
        RECT 167.000 126.200 167.300 127.800 ;
        RECT 160.600 125.800 161.000 126.200 ;
        RECT 162.200 125.800 162.600 126.200 ;
        RECT 163.000 125.800 163.400 126.200 ;
        RECT 164.600 126.100 165.000 126.200 ;
        RECT 165.400 126.100 165.800 126.200 ;
        RECT 164.600 125.800 165.800 126.100 ;
        RECT 166.200 125.800 166.600 126.200 ;
        RECT 167.000 125.800 167.400 126.200 ;
        RECT 162.200 125.200 162.500 125.800 ;
        RECT 162.200 124.800 162.600 125.200 ;
        RECT 159.800 123.800 160.200 124.200 ;
        RECT 158.200 112.100 158.600 117.900 ;
        RECT 159.800 116.200 160.100 123.800 ;
        RECT 162.200 120.800 162.600 121.200 ;
        RECT 160.600 118.100 161.000 118.200 ;
        RECT 161.400 118.100 161.800 118.200 ;
        RECT 160.600 117.800 161.800 118.100 ;
        RECT 159.800 115.800 160.200 116.200 ;
        RECT 162.200 115.200 162.500 120.800 ;
        RECT 160.600 115.100 161.000 115.200 ;
        RECT 161.400 115.100 161.800 115.200 ;
        RECT 160.600 114.800 161.800 115.100 ;
        RECT 162.200 114.800 162.600 115.200 ;
        RECT 161.400 113.800 161.800 114.200 ;
        RECT 157.400 109.800 157.800 110.200 ;
        RECT 155.800 107.800 156.200 108.200 ;
        RECT 155.000 105.800 155.400 106.200 ;
        RECT 155.800 105.900 156.200 106.300 ;
        RECT 155.000 95.200 155.300 105.800 ;
        RECT 155.800 99.200 156.100 105.900 ;
        RECT 156.600 103.100 157.000 108.900 ;
        RECT 155.800 98.800 156.200 99.200 ;
        RECT 157.400 95.200 157.700 109.800 ;
        RECT 161.400 109.200 161.700 113.800 ;
        RECT 162.200 110.200 162.500 114.800 ;
        RECT 163.000 114.200 163.300 125.800 ;
        RECT 166.200 125.200 166.500 125.800 ;
        RECT 166.200 124.800 166.600 125.200 ;
        RECT 167.000 121.200 167.300 125.800 ;
        RECT 167.000 120.800 167.400 121.200 ;
        RECT 167.000 117.800 167.400 118.200 ;
        RECT 165.400 115.800 165.800 116.200 ;
        RECT 163.000 113.800 163.400 114.200 ;
        RECT 163.000 113.100 163.400 113.200 ;
        RECT 163.800 113.100 164.200 113.200 ;
        RECT 163.000 112.800 164.200 113.100 ;
        RECT 164.600 112.800 165.000 113.200 ;
        RECT 162.200 109.800 162.600 110.200 ;
        RECT 164.600 109.200 164.900 112.800 ;
        RECT 161.400 108.800 161.800 109.200 ;
        RECT 162.200 108.800 162.600 109.200 ;
        RECT 164.600 108.800 165.000 109.200 ;
        RECT 162.200 108.100 162.500 108.800 ;
        RECT 158.200 105.100 158.600 107.900 ;
        RECT 161.400 107.800 162.500 108.100 ;
        RECT 159.000 106.800 159.400 107.200 ;
        RECT 159.000 100.200 159.300 106.800 ;
        RECT 159.800 105.800 160.200 106.200 ;
        RECT 159.800 105.200 160.100 105.800 ;
        RECT 161.400 105.200 161.700 107.800 ;
        RECT 165.400 107.200 165.700 115.800 ;
        RECT 167.000 114.200 167.300 117.800 ;
        RECT 167.000 113.800 167.400 114.200 ;
        RECT 167.800 109.200 168.100 132.800 ;
        RECT 169.400 131.800 169.800 132.200 ;
        RECT 168.600 126.800 169.000 127.200 ;
        RECT 168.600 126.200 168.900 126.800 ;
        RECT 168.600 125.800 169.000 126.200 ;
        RECT 168.600 121.800 169.000 122.200 ;
        RECT 168.600 113.100 168.900 121.800 ;
        RECT 169.400 118.200 169.700 131.800 ;
        RECT 170.200 128.200 170.500 141.800 ;
        RECT 174.200 140.800 174.600 141.200 ;
        RECT 174.200 139.200 174.500 140.800 ;
        RECT 173.400 138.800 173.800 139.200 ;
        RECT 174.200 138.800 174.600 139.200 ;
        RECT 173.400 135.200 173.700 138.800 ;
        RECT 171.000 134.800 171.400 135.200 ;
        RECT 172.600 134.800 173.000 135.200 ;
        RECT 173.400 134.800 173.800 135.200 ;
        RECT 171.000 132.200 171.300 134.800 ;
        RECT 172.600 134.200 172.900 134.800 ;
        RECT 172.600 133.800 173.000 134.200 ;
        RECT 171.000 131.800 171.400 132.200 ;
        RECT 170.200 127.800 170.600 128.200 ;
        RECT 171.000 125.100 171.400 127.900 ;
        RECT 171.800 125.800 172.200 126.200 ;
        RECT 169.400 117.800 169.800 118.200 ;
        RECT 171.000 116.800 171.400 117.200 ;
        RECT 169.400 115.800 169.800 116.200 ;
        RECT 169.400 115.200 169.700 115.800 ;
        RECT 171.000 115.200 171.300 116.800 ;
        RECT 171.800 116.100 172.100 125.800 ;
        RECT 172.600 123.100 173.000 128.900 ;
        RECT 173.400 128.200 173.700 134.800 ;
        RECT 173.400 127.800 173.800 128.200 ;
        RECT 175.000 127.200 175.300 147.800 ;
        RECT 175.800 137.200 176.100 151.800 ;
        RECT 175.800 136.800 176.200 137.200 ;
        RECT 175.800 135.800 176.200 136.200 ;
        RECT 175.800 135.200 176.100 135.800 ;
        RECT 175.800 134.800 176.200 135.200 ;
        RECT 176.600 128.200 176.900 152.800 ;
        RECT 177.400 151.200 177.700 154.800 ;
        RECT 177.400 150.800 177.800 151.200 ;
        RECT 177.400 142.100 177.800 142.200 ;
        RECT 178.200 142.100 178.600 142.200 ;
        RECT 177.400 141.800 178.600 142.100 ;
        RECT 178.200 135.800 178.600 136.200 ;
        RECT 178.200 135.200 178.500 135.800 ;
        RECT 178.200 134.800 178.600 135.200 ;
        RECT 178.200 133.800 178.600 134.200 ;
        RECT 178.200 133.200 178.500 133.800 ;
        RECT 178.200 132.800 178.600 133.200 ;
        RECT 179.800 132.800 180.200 133.200 ;
        RECT 176.600 127.800 177.000 128.200 ;
        RECT 175.000 126.800 175.400 127.200 ;
        RECT 173.400 125.900 173.800 126.300 ;
        RECT 173.400 125.200 173.700 125.900 ;
        RECT 176.600 125.800 177.000 126.200 ;
        RECT 173.400 124.800 173.800 125.200 ;
        RECT 175.000 121.800 175.400 122.200 ;
        RECT 172.600 116.100 173.000 116.200 ;
        RECT 171.800 115.800 173.000 116.100 ;
        RECT 169.400 114.800 169.800 115.200 ;
        RECT 171.000 114.800 171.400 115.200 ;
        RECT 170.200 113.800 170.600 114.200 ;
        RECT 168.600 112.800 169.700 113.100 ;
        RECT 168.600 111.800 169.000 112.200 ;
        RECT 168.600 109.200 168.900 111.800 ;
        RECT 167.800 108.800 168.200 109.200 ;
        RECT 168.600 108.800 169.000 109.200 ;
        RECT 168.600 108.100 169.000 108.200 ;
        RECT 169.400 108.100 169.700 112.800 ;
        RECT 168.600 107.800 169.700 108.100 ;
        RECT 170.200 107.200 170.500 113.800 ;
        RECT 162.200 107.100 162.600 107.200 ;
        RECT 163.000 107.100 163.400 107.200 ;
        RECT 162.200 106.800 163.400 107.100 ;
        RECT 163.800 106.800 164.200 107.200 ;
        RECT 164.600 106.800 165.000 107.200 ;
        RECT 165.400 106.800 165.800 107.200 ;
        RECT 166.200 107.100 166.600 107.200 ;
        RECT 167.000 107.100 167.400 107.200 ;
        RECT 166.200 106.800 167.400 107.100 ;
        RECT 168.600 106.800 169.000 107.200 ;
        RECT 170.200 106.800 170.600 107.200 ;
        RECT 162.200 106.100 162.600 106.200 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 162.200 105.800 163.400 106.100 ;
        RECT 159.800 104.800 160.200 105.200 ;
        RECT 161.400 104.800 161.800 105.200 ;
        RECT 163.000 102.200 163.300 105.800 ;
        RECT 163.000 101.800 163.400 102.200 ;
        RECT 163.000 100.800 163.400 101.200 ;
        RECT 159.000 99.800 159.400 100.200 ;
        RECT 159.800 98.800 160.200 99.200 ;
        RECT 159.800 95.200 160.100 98.800 ;
        RECT 160.600 96.800 161.000 97.200 ;
        RECT 160.600 96.200 160.900 96.800 ;
        RECT 160.600 95.800 161.000 96.200 ;
        RECT 163.000 95.200 163.300 100.800 ;
        RECT 163.800 95.200 164.100 106.800 ;
        RECT 164.600 106.200 164.900 106.800 ;
        RECT 164.600 105.800 165.000 106.200 ;
        RECT 165.400 105.200 165.700 106.800 ;
        RECT 166.200 105.800 166.600 106.200 ;
        RECT 165.400 104.800 165.800 105.200 ;
        RECT 165.400 101.800 165.800 102.200 ;
        RECT 155.000 94.800 155.400 95.200 ;
        RECT 157.400 94.800 157.800 95.200 ;
        RECT 158.200 94.800 158.600 95.200 ;
        RECT 159.800 94.800 160.200 95.200 ;
        RECT 162.200 94.800 162.600 95.200 ;
        RECT 163.000 94.800 163.400 95.200 ;
        RECT 163.800 95.100 164.200 95.200 ;
        RECT 164.600 95.100 165.000 95.200 ;
        RECT 163.800 94.800 165.000 95.100 ;
        RECT 158.200 94.200 158.500 94.800 ;
        RECT 162.200 94.200 162.500 94.800 ;
        RECT 158.200 93.800 158.600 94.200 ;
        RECT 162.200 93.800 162.600 94.200 ;
        RECT 152.600 91.800 153.000 92.200 ;
        RECT 152.600 91.200 152.900 91.800 ;
        RECT 152.600 90.800 153.000 91.200 ;
        RECT 151.000 90.100 151.400 90.200 ;
        RECT 150.200 89.800 151.400 90.100 ;
        RECT 163.000 89.200 163.300 94.800 ;
        RECT 164.600 91.800 165.000 92.200 ;
        RECT 140.600 87.800 141.000 88.200 ;
        RECT 144.600 87.800 145.000 88.200 ;
        RECT 134.200 85.800 134.600 86.200 ;
        RECT 137.400 85.800 137.800 86.200 ;
        RECT 131.800 81.800 132.200 82.200 ;
        RECT 132.600 82.100 133.000 82.200 ;
        RECT 133.400 82.100 133.800 82.200 ;
        RECT 132.600 81.800 133.800 82.100 ;
        RECT 127.800 80.800 128.200 81.200 ;
        RECT 128.600 76.800 129.000 77.200 ;
        RECT 131.000 76.800 131.400 77.200 ;
        RECT 128.600 75.200 128.900 76.800 ;
        RECT 125.400 74.800 125.800 75.200 ;
        RECT 126.200 75.100 126.600 75.200 ;
        RECT 127.000 75.100 127.400 75.200 ;
        RECT 126.200 74.800 127.400 75.100 ;
        RECT 128.600 74.800 129.000 75.200 ;
        RECT 129.400 74.800 129.800 75.200 ;
        RECT 124.600 73.800 125.000 74.200 ;
        RECT 123.800 70.800 124.200 71.200 ;
        RECT 121.400 67.800 121.800 68.200 ;
        RECT 121.400 67.200 121.700 67.800 ;
        RECT 121.400 66.800 121.800 67.200 ;
        RECT 123.000 66.800 123.400 67.200 ;
        RECT 123.800 66.800 124.200 67.200 ;
        RECT 123.000 66.200 123.300 66.800 ;
        RECT 123.800 66.200 124.100 66.800 ;
        RECT 118.200 66.100 118.600 66.200 ;
        RECT 119.000 66.100 119.400 66.200 ;
        RECT 118.200 65.800 119.400 66.100 ;
        RECT 119.800 65.800 120.200 66.200 ;
        RECT 120.600 65.800 121.000 66.200 ;
        RECT 123.000 65.800 123.400 66.200 ;
        RECT 123.800 65.800 124.200 66.200 ;
        RECT 119.800 65.200 120.100 65.800 ;
        RECT 119.800 64.800 120.200 65.200 ;
        RECT 117.400 58.800 117.800 59.200 ;
        RECT 118.200 58.800 118.600 59.200 ;
        RECT 119.000 58.800 119.400 59.200 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 114.200 55.100 114.600 55.200 ;
        RECT 115.000 55.100 115.400 55.200 ;
        RECT 114.200 54.800 115.400 55.100 ;
        RECT 115.800 54.800 116.200 55.200 ;
        RECT 111.800 54.200 112.100 54.800 ;
        RECT 118.200 54.200 118.500 58.800 ;
        RECT 119.000 58.200 119.300 58.800 ;
        RECT 119.000 57.800 119.400 58.200 ;
        RECT 120.600 55.200 120.900 65.800 ;
        RECT 124.600 65.100 125.000 67.900 ;
        RECT 121.400 61.800 121.800 62.200 ;
        RECT 121.400 59.200 121.700 61.800 ;
        RECT 123.800 59.800 124.200 60.200 ;
        RECT 121.400 58.800 121.800 59.200 ;
        RECT 123.800 55.200 124.100 59.800 ;
        RECT 119.000 54.800 119.400 55.200 ;
        RECT 120.600 54.800 121.000 55.200 ;
        RECT 123.800 54.800 124.200 55.200 ;
        RECT 111.800 53.800 112.200 54.200 ;
        RECT 118.200 53.800 118.600 54.200 ;
        RECT 110.200 52.800 110.600 53.200 ;
        RECT 116.600 52.800 117.000 53.200 ;
        RECT 110.200 51.800 110.600 52.200 ;
        RECT 107.800 49.800 108.200 50.200 ;
        RECT 107.800 48.200 108.100 49.800 ;
        RECT 108.600 49.100 109.000 49.200 ;
        RECT 109.400 49.100 109.800 49.200 ;
        RECT 108.600 48.800 109.800 49.100 ;
        RECT 104.600 47.800 105.000 48.200 ;
        RECT 107.800 47.800 108.200 48.200 ;
        RECT 108.600 47.800 109.000 48.200 ;
        RECT 104.600 46.800 105.000 47.200 ;
        RECT 106.200 46.800 106.600 47.200 ;
        RECT 101.400 45.800 101.800 46.200 ;
        RECT 102.200 46.100 102.600 46.200 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 102.200 45.800 103.400 46.100 ;
        RECT 100.600 42.800 101.000 43.200 ;
        RECT 101.400 40.200 101.700 45.800 ;
        RECT 104.600 43.200 104.900 46.800 ;
        RECT 105.400 45.800 105.800 46.200 ;
        RECT 104.600 42.800 105.000 43.200 ;
        RECT 101.400 39.800 101.800 40.200 ;
        RECT 103.000 39.100 103.400 39.200 ;
        RECT 103.800 39.100 104.200 39.200 ;
        RECT 103.000 38.800 104.200 39.100 ;
        RECT 100.600 35.800 101.000 36.200 ;
        RECT 100.600 29.200 100.900 35.800 ;
        RECT 101.400 32.100 101.800 37.900 ;
        RECT 104.600 36.800 105.000 37.200 ;
        RECT 104.600 33.200 104.900 36.800 ;
        RECT 103.800 33.100 104.200 33.200 ;
        RECT 104.600 33.100 105.000 33.200 ;
        RECT 103.800 32.800 105.000 33.100 ;
        RECT 100.600 28.800 101.000 29.200 ;
        RECT 100.600 26.200 100.900 28.800 ;
        RECT 105.400 28.200 105.700 45.800 ;
        RECT 106.200 38.200 106.500 46.800 ;
        RECT 107.000 41.800 107.400 42.200 ;
        RECT 106.200 37.800 106.600 38.200 ;
        RECT 107.000 35.200 107.300 41.800 ;
        RECT 106.200 34.800 106.600 35.200 ;
        RECT 107.000 34.800 107.400 35.200 ;
        RECT 106.200 34.200 106.500 34.800 ;
        RECT 108.600 34.200 108.900 47.800 ;
        RECT 109.400 45.100 109.800 47.900 ;
        RECT 110.200 47.200 110.500 51.800 ;
        RECT 116.600 51.200 116.900 52.800 ;
        RECT 116.600 50.800 117.000 51.200 ;
        RECT 118.200 49.800 118.600 50.200 ;
        RECT 118.200 49.200 118.500 49.800 ;
        RECT 119.000 49.200 119.300 54.800 ;
        RECT 123.800 54.100 124.200 54.200 ;
        RECT 124.600 54.100 125.000 54.200 ;
        RECT 123.800 53.800 125.000 54.100 ;
        RECT 122.200 49.800 122.600 50.200 ;
        RECT 110.200 46.800 110.600 47.200 ;
        RECT 111.000 43.100 111.400 48.900 ;
        RECT 112.600 46.800 113.000 47.200 ;
        RECT 112.600 46.200 112.900 46.800 ;
        RECT 112.600 45.800 113.000 46.200 ;
        RECT 115.800 43.100 116.200 48.900 ;
        RECT 118.200 48.800 118.600 49.200 ;
        RECT 119.000 48.800 119.400 49.200 ;
        RECT 121.400 48.800 121.800 49.200 ;
        RECT 120.600 47.800 121.000 48.200 ;
        RECT 120.600 46.200 120.900 47.800 ;
        RECT 121.400 47.200 121.700 48.800 ;
        RECT 122.200 48.200 122.500 49.800 ;
        RECT 123.800 48.800 124.200 49.200 ;
        RECT 122.200 47.800 122.600 48.200 ;
        RECT 123.800 47.200 124.100 48.800 ;
        RECT 121.400 46.800 121.800 47.200 ;
        RECT 123.800 46.800 124.200 47.200 ;
        RECT 120.600 45.800 121.000 46.200 ;
        RECT 122.200 45.800 122.600 46.200 ;
        RECT 123.800 46.100 124.200 46.200 ;
        RECT 124.600 46.100 125.000 46.200 ;
        RECT 123.800 45.800 125.000 46.100 ;
        RECT 116.600 44.800 117.000 45.200 ;
        RECT 118.200 45.100 118.600 45.200 ;
        RECT 119.000 45.100 119.400 45.200 ;
        RECT 118.200 44.800 119.400 45.100 ;
        RECT 120.600 44.800 121.000 45.200 ;
        RECT 109.400 37.100 109.800 37.200 ;
        RECT 110.200 37.100 110.600 37.200 ;
        RECT 109.400 36.800 110.600 37.100 ;
        RECT 109.400 34.800 109.800 35.200 ;
        RECT 106.200 33.800 106.600 34.200 ;
        RECT 108.600 33.800 109.000 34.200 ;
        RECT 107.800 32.800 108.200 33.200 ;
        RECT 107.800 32.200 108.100 32.800 ;
        RECT 107.800 31.800 108.200 32.200 ;
        RECT 107.800 30.800 108.200 31.200 ;
        RECT 105.400 27.800 105.800 28.200 ;
        RECT 103.800 26.800 104.200 27.200 ;
        RECT 103.800 26.200 104.100 26.800 ;
        RECT 97.400 26.100 97.800 26.200 ;
        RECT 98.200 26.100 98.600 26.200 ;
        RECT 97.400 25.800 98.600 26.100 ;
        RECT 99.800 25.800 100.200 26.200 ;
        RECT 100.600 25.800 101.000 26.200 ;
        RECT 103.800 25.800 104.200 26.200 ;
        RECT 99.800 21.200 100.100 25.800 ;
        RECT 96.600 20.800 97.000 21.200 ;
        RECT 99.800 20.800 100.200 21.200 ;
        RECT 91.000 18.800 91.400 19.200 ;
        RECT 87.800 16.800 88.200 17.200 ;
        RECT 87.800 14.200 88.100 16.800 ;
        RECT 87.800 13.800 88.200 14.200 ;
        RECT 88.600 13.100 89.000 15.900 ;
        RECT 91.000 13.200 91.300 18.800 ;
        RECT 95.800 15.800 96.200 16.200 ;
        RECT 95.800 15.200 96.100 15.800 ;
        RECT 96.600 15.200 96.900 20.800 ;
        RECT 97.400 19.100 97.800 19.200 ;
        RECT 98.200 19.100 98.600 19.200 ;
        RECT 97.400 18.800 98.600 19.100 ;
        RECT 107.000 18.800 107.400 19.200 ;
        RECT 92.600 14.800 93.000 15.200 ;
        RECT 95.000 14.800 95.400 15.200 ;
        RECT 95.800 14.800 96.200 15.200 ;
        RECT 96.600 14.800 97.000 15.200 ;
        RECT 92.600 14.200 92.900 14.800 ;
        RECT 92.600 13.800 93.000 14.200 ;
        RECT 91.000 12.800 91.400 13.200 ;
        RECT 95.000 9.200 95.300 14.800 ;
        RECT 99.800 12.100 100.200 17.900 ;
        RECT 100.600 16.800 101.000 17.200 ;
        RECT 100.600 15.200 100.900 16.800 ;
        RECT 103.800 15.800 104.200 16.200 ;
        RECT 100.600 14.800 101.000 15.200 ;
        RECT 103.800 15.100 104.100 15.800 ;
        RECT 103.800 14.700 104.200 15.100 ;
        RECT 104.600 12.100 105.000 17.900 ;
        RECT 106.200 13.100 106.600 15.900 ;
        RECT 107.000 13.200 107.300 18.800 ;
        RECT 107.000 12.800 107.400 13.200 ;
        RECT 107.800 12.100 108.100 30.800 ;
        RECT 108.600 23.100 109.000 28.900 ;
        RECT 109.400 15.200 109.700 34.800 ;
        RECT 112.600 32.100 113.000 37.900 ;
        RECT 114.200 34.800 114.600 35.200 ;
        RECT 114.200 33.200 114.500 34.800 ;
        RECT 115.800 33.800 116.200 34.200 ;
        RECT 114.200 32.800 114.600 33.200 ;
        RECT 111.000 26.100 111.400 26.200 ;
        RECT 111.800 26.100 112.200 26.200 ;
        RECT 111.000 25.800 112.200 26.100 ;
        RECT 113.400 23.100 113.800 28.900 ;
        RECT 114.200 26.800 114.600 27.200 ;
        RECT 114.200 26.200 114.500 26.800 ;
        RECT 114.200 25.800 114.600 26.200 ;
        RECT 115.000 25.100 115.400 27.900 ;
        RECT 115.800 26.200 116.100 33.800 ;
        RECT 116.600 29.200 116.900 44.800 ;
        RECT 120.600 39.200 120.900 44.800 ;
        RECT 120.600 38.800 121.000 39.200 ;
        RECT 117.400 32.100 117.800 37.900 ;
        RECT 122.200 36.200 122.500 45.800 ;
        RECT 125.400 39.200 125.700 74.800 ;
        RECT 129.400 74.200 129.700 74.800 ;
        RECT 129.400 73.800 129.800 74.200 ;
        RECT 131.000 73.200 131.300 76.800 ;
        RECT 131.000 72.800 131.400 73.200 ;
        RECT 127.000 69.800 127.400 70.200 ;
        RECT 126.200 63.100 126.600 68.900 ;
        RECT 127.000 68.200 127.300 69.800 ;
        RECT 127.000 67.800 127.400 68.200 ;
        RECT 127.000 65.900 127.400 66.300 ;
        RECT 127.000 65.200 127.300 65.900 ;
        RECT 127.000 64.800 127.400 65.200 ;
        RECT 131.000 63.100 131.400 68.900 ;
        RECT 131.000 60.800 131.400 61.200 ;
        RECT 126.200 52.800 126.600 53.200 ;
        RECT 126.200 49.200 126.500 52.800 ;
        RECT 127.000 52.100 127.400 52.200 ;
        RECT 127.800 52.100 128.200 52.200 ;
        RECT 129.400 52.100 129.800 57.900 ;
        RECT 130.200 54.800 130.600 55.200 ;
        RECT 127.000 51.800 128.200 52.100 ;
        RECT 126.200 48.800 126.600 49.200 ;
        RECT 127.000 47.100 127.400 47.200 ;
        RECT 127.800 47.100 128.200 47.200 ;
        RECT 127.000 46.800 128.200 47.100 ;
        RECT 130.200 46.200 130.500 54.800 ;
        RECT 131.000 47.200 131.300 60.800 ;
        RECT 131.800 48.200 132.100 81.800 ;
        RECT 133.400 80.800 133.800 81.200 ;
        RECT 133.400 79.200 133.700 80.800 ;
        RECT 133.400 78.800 133.800 79.200 ;
        RECT 132.600 75.800 133.000 76.200 ;
        RECT 132.600 75.200 132.900 75.800 ;
        RECT 132.600 74.800 133.000 75.200 ;
        RECT 132.600 73.200 132.900 74.800 ;
        RECT 132.600 72.800 133.000 73.200 ;
        RECT 134.200 72.200 134.500 85.800 ;
        RECT 137.400 85.200 137.700 85.800 ;
        RECT 137.400 84.800 137.800 85.200 ;
        RECT 145.400 82.100 145.800 88.900 ;
        RECT 146.200 82.100 146.600 88.900 ;
        RECT 147.000 83.100 147.400 88.900 ;
        RECT 147.800 88.800 148.200 89.200 ;
        RECT 160.600 89.100 161.000 89.200 ;
        RECT 161.400 89.100 161.800 89.200 ;
        RECT 147.800 87.200 148.100 88.800 ;
        RECT 147.800 86.800 148.200 87.200 ;
        RECT 148.600 83.100 149.000 88.900 ;
        RECT 149.400 87.800 149.800 88.200 ;
        RECT 149.400 87.200 149.700 87.800 ;
        RECT 149.400 86.800 149.800 87.200 ;
        RECT 150.200 83.100 150.600 88.900 ;
        RECT 151.000 82.100 151.400 88.900 ;
        RECT 151.800 82.100 152.200 88.900 ;
        RECT 152.600 82.100 153.000 88.900 ;
        RECT 160.600 88.800 161.800 89.100 ;
        RECT 163.000 88.800 163.400 89.200 ;
        RECT 157.400 88.100 157.800 88.200 ;
        RECT 158.200 88.100 158.600 88.200 ;
        RECT 157.400 87.800 158.600 88.100 ;
        RECT 163.800 87.800 164.200 88.200 ;
        RECT 163.800 87.200 164.100 87.800 ;
        RECT 164.600 87.200 164.900 91.800 ;
        RECT 159.000 87.100 159.400 87.200 ;
        RECT 159.800 87.100 160.200 87.200 ;
        RECT 159.000 86.800 160.200 87.100 ;
        RECT 163.800 86.800 164.200 87.200 ;
        RECT 164.600 86.800 165.000 87.200 ;
        RECT 165.400 86.200 165.700 101.800 ;
        RECT 166.200 92.200 166.500 105.800 ;
        RECT 167.000 104.800 167.400 105.200 ;
        RECT 166.200 91.800 166.600 92.200 ;
        RECT 167.000 91.100 167.300 104.800 ;
        RECT 167.800 92.100 168.200 97.900 ;
        RECT 167.000 90.800 168.100 91.100 ;
        RECT 167.000 88.800 167.400 89.200 ;
        RECT 167.000 88.200 167.300 88.800 ;
        RECT 167.000 87.800 167.400 88.200 ;
        RECT 167.800 87.200 168.100 90.800 ;
        RECT 168.600 87.200 168.900 106.800 ;
        RECT 169.400 106.100 169.800 106.200 ;
        RECT 170.200 106.100 170.600 106.200 ;
        RECT 169.400 105.800 170.600 106.100 ;
        RECT 171.000 95.800 171.400 96.200 ;
        RECT 171.000 95.200 171.300 95.800 ;
        RECT 171.000 94.800 171.400 95.200 ;
        RECT 171.000 87.800 171.400 88.200 ;
        RECT 167.800 86.800 168.200 87.200 ;
        RECT 168.600 86.800 169.000 87.200 ;
        RECT 159.000 86.100 159.400 86.200 ;
        RECT 159.000 85.800 160.100 86.100 ;
        RECT 135.800 79.800 136.200 80.200 ;
        RECT 135.000 75.800 135.400 76.200 ;
        RECT 135.000 75.200 135.300 75.800 ;
        RECT 135.800 75.200 136.100 79.800 ;
        RECT 139.000 77.800 139.400 78.200 ;
        RECT 137.400 77.100 137.800 77.200 ;
        RECT 138.200 77.100 138.600 77.200 ;
        RECT 137.400 76.800 138.600 77.100 ;
        RECT 135.000 74.800 135.400 75.200 ;
        RECT 135.800 74.800 136.200 75.200 ;
        RECT 137.400 74.800 137.800 75.200 ;
        RECT 134.200 71.800 134.600 72.200 ;
        RECT 135.800 67.800 136.200 68.200 ;
        RECT 135.800 67.200 136.100 67.800 ;
        RECT 134.200 66.800 134.600 67.200 ;
        RECT 135.800 66.800 136.200 67.200 ;
        RECT 134.200 66.200 134.500 66.800 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 135.000 66.100 135.400 66.200 ;
        RECT 134.200 65.800 135.400 66.100 ;
        RECT 135.800 66.100 136.200 66.200 ;
        RECT 136.600 66.100 137.000 66.200 ;
        RECT 135.800 65.800 137.000 66.100 ;
        RECT 137.400 63.200 137.700 74.800 ;
        RECT 138.200 70.800 138.600 71.200 ;
        RECT 138.200 66.200 138.500 70.800 ;
        RECT 139.000 67.200 139.300 77.800 ;
        RECT 140.600 72.100 141.000 77.900 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 143.000 75.100 143.400 75.200 ;
        RECT 143.800 75.100 144.200 75.200 ;
        RECT 143.000 74.800 144.200 75.100 ;
        RECT 141.400 68.800 141.800 69.200 ;
        RECT 141.400 67.200 141.700 68.800 ;
        RECT 139.000 66.800 139.400 67.200 ;
        RECT 141.400 66.800 141.800 67.200 ;
        RECT 142.200 66.200 142.500 74.800 ;
        RECT 144.600 72.800 145.000 73.200 ;
        RECT 144.600 71.100 144.900 72.800 ;
        RECT 145.400 72.100 145.800 77.900 ;
        RECT 147.000 73.100 147.400 75.900 ;
        RECT 147.000 71.800 147.400 72.200 ;
        RECT 151.800 72.100 152.200 78.900 ;
        RECT 152.600 72.100 153.000 78.900 ;
        RECT 153.400 72.100 153.800 77.900 ;
        RECT 154.200 73.800 154.600 74.200 ;
        RECT 144.600 70.800 145.700 71.100 ;
        RECT 143.800 67.800 144.200 68.200 ;
        RECT 143.800 66.200 144.100 67.800 ;
        RECT 144.600 66.800 145.000 67.200 ;
        RECT 138.200 65.800 138.600 66.200 ;
        RECT 142.200 65.800 142.600 66.200 ;
        RECT 143.800 65.800 144.200 66.200 ;
        RECT 137.400 62.800 137.800 63.200 ;
        RECT 136.600 61.800 137.000 62.200 ;
        RECT 138.200 62.100 138.500 65.800 ;
        RECT 137.400 61.800 138.500 62.100 ;
        RECT 136.600 60.200 136.900 61.800 ;
        RECT 136.600 59.800 137.000 60.200 ;
        RECT 132.600 57.800 133.000 58.200 ;
        RECT 132.600 49.200 132.900 57.800 ;
        RECT 133.400 55.800 133.800 56.200 ;
        RECT 133.400 55.100 133.700 55.800 ;
        RECT 133.400 54.700 133.800 55.100 ;
        RECT 134.200 52.100 134.600 57.900 ;
        RECT 135.000 54.800 135.400 55.200 ;
        RECT 135.000 54.200 135.300 54.800 ;
        RECT 135.000 53.800 135.400 54.200 ;
        RECT 135.800 53.100 136.200 55.900 ;
        RECT 136.600 52.800 137.000 53.200 ;
        RECT 136.600 52.200 136.900 52.800 ;
        RECT 136.600 51.800 137.000 52.200 ;
        RECT 132.600 48.800 133.000 49.200 ;
        RECT 131.800 47.800 132.200 48.200 ;
        RECT 136.600 47.800 137.000 48.200 ;
        RECT 131.000 46.800 131.400 47.200 ;
        RECT 133.400 46.800 133.800 47.200 ;
        RECT 134.200 46.800 134.600 47.200 ;
        RECT 131.000 46.200 131.300 46.800 ;
        RECT 133.400 46.200 133.700 46.800 ;
        RECT 134.200 46.200 134.500 46.800 ;
        RECT 136.600 46.200 136.900 47.800 ;
        RECT 127.000 46.100 127.400 46.200 ;
        RECT 127.800 46.100 128.200 46.200 ;
        RECT 127.000 45.800 128.200 46.100 ;
        RECT 130.200 45.800 130.600 46.200 ;
        RECT 131.000 45.800 131.400 46.200 ;
        RECT 133.400 45.800 133.800 46.200 ;
        RECT 134.200 45.800 134.600 46.200 ;
        RECT 136.600 45.800 137.000 46.200 ;
        RECT 126.200 44.800 126.600 45.200 ;
        RECT 125.400 38.800 125.800 39.200 ;
        RECT 119.000 33.100 119.400 35.900 ;
        RECT 122.200 35.800 122.600 36.200 ;
        RECT 122.200 35.200 122.500 35.800 ;
        RECT 119.800 35.100 120.200 35.200 ;
        RECT 120.600 35.100 121.000 35.200 ;
        RECT 119.800 34.800 121.000 35.100 ;
        RECT 122.200 34.800 122.600 35.200 ;
        RECT 119.800 34.100 120.200 34.200 ;
        RECT 120.600 34.100 121.000 34.200 ;
        RECT 119.800 33.800 121.000 34.100 ;
        RECT 123.800 33.800 124.200 34.200 ;
        RECT 122.200 33.100 122.600 33.200 ;
        RECT 123.000 33.100 123.400 33.200 ;
        RECT 122.200 32.800 123.400 33.100 ;
        RECT 123.800 31.200 124.100 33.800 ;
        RECT 125.400 31.800 125.800 32.200 ;
        RECT 125.400 31.200 125.700 31.800 ;
        RECT 123.800 30.800 124.200 31.200 ;
        RECT 125.400 30.800 125.800 31.200 ;
        RECT 126.200 30.100 126.500 44.800 ;
        RECT 125.400 29.800 126.500 30.100 ;
        RECT 127.000 33.800 127.400 34.200 ;
        RECT 127.000 32.200 127.300 33.800 ;
        RECT 127.000 31.800 127.400 32.200 ;
        RECT 125.400 29.200 125.700 29.800 ;
        RECT 116.600 28.800 117.000 29.200 ;
        RECT 119.000 28.800 119.400 29.200 ;
        RECT 125.400 28.800 125.800 29.200 ;
        RECT 117.400 26.800 117.800 27.200 ;
        RECT 115.800 25.800 116.200 26.200 ;
        RECT 115.800 25.100 116.200 25.200 ;
        RECT 116.600 25.100 117.000 25.200 ;
        RECT 115.800 24.800 117.000 25.100 ;
        RECT 112.600 20.800 113.000 21.200 ;
        RECT 111.800 19.800 112.200 20.200 ;
        RECT 110.200 16.800 110.600 17.200 ;
        RECT 110.200 16.200 110.500 16.800 ;
        RECT 110.200 15.800 110.600 16.200 ;
        RECT 111.800 15.200 112.100 19.800 ;
        RECT 112.600 15.200 112.900 20.800 ;
        RECT 117.400 16.200 117.700 26.800 ;
        RECT 119.000 26.200 119.300 28.800 ;
        RECT 123.800 28.100 124.200 28.200 ;
        RECT 124.600 28.100 125.000 28.200 ;
        RECT 123.800 27.800 125.000 28.100 ;
        RECT 126.200 27.800 126.600 28.200 ;
        RECT 126.200 27.200 126.500 27.800 ;
        RECT 121.400 27.100 121.800 27.200 ;
        RECT 122.200 27.100 122.600 27.200 ;
        RECT 121.400 26.800 122.600 27.100 ;
        RECT 126.200 26.800 126.600 27.200 ;
        RECT 127.000 26.200 127.300 31.800 ;
        RECT 130.200 29.200 130.500 45.800 ;
        RECT 136.600 43.800 137.000 44.200 ;
        RECT 135.800 41.800 136.200 42.200 ;
        RECT 133.400 33.100 133.800 35.900 ;
        RECT 134.200 33.800 134.600 34.200 ;
        RECT 134.200 33.200 134.500 33.800 ;
        RECT 134.200 32.800 134.600 33.200 ;
        RECT 135.000 32.100 135.400 37.900 ;
        RECT 135.800 35.100 136.100 41.800 ;
        RECT 135.800 34.700 136.200 35.100 ;
        RECT 136.600 29.200 136.900 43.800 ;
        RECT 137.400 32.200 137.700 61.800 ;
        RECT 142.200 58.200 142.500 65.800 ;
        RECT 143.000 65.100 143.400 65.200 ;
        RECT 143.800 65.100 144.200 65.200 ;
        RECT 143.000 64.800 144.200 65.100 ;
        RECT 144.600 62.200 144.900 66.800 ;
        RECT 143.000 61.800 143.400 62.200 ;
        RECT 144.600 61.800 145.000 62.200 ;
        RECT 142.200 57.800 142.600 58.200 ;
        RECT 143.000 56.200 143.300 61.800 ;
        RECT 138.200 56.100 138.600 56.200 ;
        RECT 139.000 56.100 139.400 56.200 ;
        RECT 138.200 55.800 139.400 56.100 ;
        RECT 143.000 55.800 143.400 56.200 ;
        RECT 143.800 55.800 144.200 56.200 ;
        RECT 143.000 55.200 143.300 55.800 ;
        RECT 143.800 55.200 144.100 55.800 ;
        RECT 138.200 54.800 138.600 55.200 ;
        RECT 140.600 55.100 141.000 55.200 ;
        RECT 141.400 55.100 141.800 55.200 ;
        RECT 140.600 54.800 141.800 55.100 ;
        RECT 143.000 54.800 143.400 55.200 ;
        RECT 143.800 54.800 144.200 55.200 ;
        RECT 138.200 54.200 138.500 54.800 ;
        RECT 138.200 53.800 138.600 54.200 ;
        RECT 142.200 53.800 142.600 54.200 ;
        RECT 142.200 49.200 142.500 53.800 ;
        RECT 143.800 51.200 144.100 54.800 ;
        RECT 144.600 53.100 145.000 55.900 ;
        RECT 145.400 54.200 145.700 70.800 ;
        RECT 147.000 69.200 147.300 71.800 ;
        RECT 154.200 71.100 154.500 73.800 ;
        RECT 155.000 72.100 155.400 77.900 ;
        RECT 155.800 72.800 156.200 73.200 ;
        RECT 155.800 72.200 156.100 72.800 ;
        RECT 155.800 71.800 156.200 72.200 ;
        RECT 156.600 72.100 157.000 77.900 ;
        RECT 157.400 72.100 157.800 78.900 ;
        RECT 158.200 72.100 158.600 78.900 ;
        RECT 159.000 72.100 159.400 78.900 ;
        RECT 153.400 70.800 154.500 71.100 ;
        RECT 153.400 69.200 153.700 70.800 ;
        RECT 155.000 69.800 155.400 70.200 ;
        RECT 147.000 68.800 147.400 69.200 ;
        RECT 153.400 68.800 153.800 69.200 ;
        RECT 154.200 68.800 154.600 69.200 ;
        RECT 154.200 68.200 154.500 68.800 ;
        RECT 146.200 67.800 146.600 68.200 ;
        RECT 151.800 67.800 153.700 68.100 ;
        RECT 154.200 67.800 154.600 68.200 ;
        RECT 146.200 64.200 146.500 67.800 ;
        RECT 151.800 67.200 152.100 67.800 ;
        RECT 147.800 67.100 148.200 67.200 ;
        RECT 150.200 67.100 150.600 67.200 ;
        RECT 147.800 66.800 150.600 67.100 ;
        RECT 151.800 66.800 152.200 67.200 ;
        RECT 152.600 66.800 153.000 67.200 ;
        RECT 153.400 67.100 153.700 67.800 ;
        RECT 154.200 67.100 154.600 67.200 ;
        RECT 153.400 66.800 154.600 67.100 ;
        RECT 147.800 65.800 148.200 66.200 ;
        RECT 151.800 65.800 152.200 66.200 ;
        RECT 147.800 65.200 148.100 65.800 ;
        RECT 147.800 64.800 148.200 65.200 ;
        RECT 146.200 63.800 146.600 64.200 ;
        RECT 151.800 60.200 152.100 65.800 ;
        RECT 152.600 65.200 152.900 66.800 ;
        RECT 155.000 65.200 155.300 69.800 ;
        RECT 157.400 66.800 157.800 67.200 ;
        RECT 152.600 64.800 153.000 65.200 ;
        RECT 155.000 64.800 155.400 65.200 ;
        RECT 154.200 62.800 154.600 63.200 ;
        RECT 151.800 59.800 152.200 60.200 ;
        RECT 145.400 53.800 145.800 54.200 ;
        RECT 145.400 53.200 145.700 53.800 ;
        RECT 145.400 52.800 145.800 53.200 ;
        RECT 146.200 52.100 146.600 57.900 ;
        RECT 147.800 57.800 148.200 58.200 ;
        RECT 147.800 55.200 148.100 57.800 ;
        RECT 149.400 56.800 149.800 57.200 ;
        RECT 147.800 54.800 148.200 55.200 ;
        RECT 143.800 50.800 144.200 51.200 ;
        RECT 142.200 48.800 142.600 49.200 ;
        RECT 140.600 47.800 141.000 48.200 ;
        RECT 146.200 47.800 146.600 48.200 ;
        RECT 140.600 39.200 140.900 47.800 ;
        RECT 146.200 39.200 146.500 47.800 ;
        RECT 149.400 46.200 149.700 56.800 ;
        RECT 150.200 53.800 150.600 54.200 ;
        RECT 150.200 46.200 150.500 53.800 ;
        RECT 151.000 52.100 151.400 57.900 ;
        RECT 154.200 55.200 154.500 62.800 ;
        RECT 157.400 59.200 157.700 66.800 ;
        RECT 158.200 65.800 158.600 66.200 ;
        RECT 157.400 58.800 157.800 59.200 ;
        RECT 157.400 56.800 157.800 57.200 ;
        RECT 157.400 55.200 157.700 56.800 ;
        RECT 154.200 54.800 154.600 55.200 ;
        RECT 155.000 55.100 155.400 55.200 ;
        RECT 155.800 55.100 156.200 55.200 ;
        RECT 155.000 54.800 156.200 55.100 ;
        RECT 157.400 54.800 157.800 55.200 ;
        RECT 154.200 52.200 154.500 54.800 ;
        RECT 155.800 53.800 156.200 54.200 ;
        RECT 153.400 51.800 153.800 52.200 ;
        RECT 154.200 51.800 154.600 52.200 ;
        RECT 153.400 51.200 153.700 51.800 ;
        RECT 153.400 50.800 153.800 51.200 ;
        RECT 155.000 50.800 155.400 51.200 ;
        RECT 153.400 46.800 153.800 47.200 ;
        RECT 148.600 45.800 149.000 46.200 ;
        RECT 149.400 45.800 149.800 46.200 ;
        RECT 150.200 45.800 150.600 46.200 ;
        RECT 151.800 45.800 152.200 46.200 ;
        RECT 148.600 42.200 148.900 45.800 ;
        RECT 148.600 41.800 149.000 42.200 ;
        RECT 140.600 38.800 141.000 39.200 ;
        RECT 141.400 39.100 141.800 39.200 ;
        RECT 142.200 39.100 142.600 39.200 ;
        RECT 141.400 38.800 142.600 39.100 ;
        RECT 146.200 38.800 146.600 39.200 ;
        RECT 149.400 39.100 149.700 45.800 ;
        RECT 148.600 38.800 149.700 39.100 ;
        RECT 137.400 31.800 137.800 32.200 ;
        RECT 139.000 31.800 139.400 32.200 ;
        RECT 139.800 32.100 140.200 37.900 ;
        RECT 143.000 36.100 143.400 36.200 ;
        RECT 142.200 35.800 143.400 36.100 ;
        RECT 118.200 25.800 118.600 26.200 ;
        RECT 119.000 25.800 119.400 26.200 ;
        RECT 127.000 25.800 127.400 26.200 ;
        RECT 118.200 21.200 118.500 25.800 ;
        RECT 118.200 20.800 118.600 21.200 ;
        RECT 113.400 16.100 113.800 16.200 ;
        RECT 114.200 16.100 114.600 16.200 ;
        RECT 113.400 15.800 114.600 16.100 ;
        RECT 115.800 15.800 116.200 16.200 ;
        RECT 117.400 15.800 117.800 16.200 ;
        RECT 115.800 15.200 116.100 15.800 ;
        RECT 109.400 14.800 109.800 15.200 ;
        RECT 111.800 14.800 112.200 15.200 ;
        RECT 112.600 14.800 113.000 15.200 ;
        RECT 115.000 14.800 115.400 15.200 ;
        RECT 115.800 14.800 116.200 15.200 ;
        RECT 117.400 15.100 117.800 15.200 ;
        RECT 118.200 15.100 118.600 15.200 ;
        RECT 119.000 15.100 119.300 25.800 ;
        RECT 123.800 25.100 124.200 25.200 ;
        RECT 124.600 25.100 125.000 25.200 ;
        RECT 123.800 24.800 125.000 25.100 ;
        RECT 121.400 20.800 121.800 21.200 ;
        RECT 121.400 15.200 121.700 20.800 ;
        RECT 122.200 15.800 122.600 16.200 ;
        RECT 122.200 15.200 122.500 15.800 ;
        RECT 117.400 14.800 119.300 15.100 ;
        RECT 119.800 15.100 120.200 15.200 ;
        RECT 120.600 15.100 121.000 15.200 ;
        RECT 119.800 14.800 121.000 15.100 ;
        RECT 121.400 14.800 121.800 15.200 ;
        RECT 122.200 14.800 122.600 15.200 ;
        RECT 123.800 15.100 124.200 15.200 ;
        RECT 124.600 15.100 125.000 15.200 ;
        RECT 123.800 14.800 125.000 15.100 ;
        RECT 115.000 14.200 115.300 14.800 ;
        RECT 115.000 13.800 115.400 14.200 ;
        RECT 113.400 12.800 113.800 13.200 ;
        RECT 117.400 12.800 117.800 13.200 ;
        RECT 119.000 13.100 119.400 13.200 ;
        RECT 119.800 13.100 120.200 13.200 ;
        RECT 126.200 13.100 126.600 15.900 ;
        RECT 127.000 14.200 127.300 25.800 ;
        RECT 129.400 23.100 129.800 28.900 ;
        RECT 130.200 28.800 130.600 29.200 ;
        RECT 132.600 26.800 133.000 27.200 ;
        RECT 132.600 26.200 132.900 26.800 ;
        RECT 130.200 25.800 130.600 26.200 ;
        RECT 132.600 25.800 133.000 26.200 ;
        RECT 130.200 25.200 130.500 25.800 ;
        RECT 130.200 24.800 130.600 25.200 ;
        RECT 134.200 23.100 134.600 28.900 ;
        RECT 136.600 28.800 137.000 29.200 ;
        RECT 135.800 25.100 136.200 27.900 ;
        RECT 139.000 27.200 139.300 31.800 ;
        RECT 142.200 29.200 142.500 35.800 ;
        RECT 146.200 34.800 146.600 35.200 ;
        RECT 143.000 30.800 143.400 31.200 ;
        RECT 142.200 28.800 142.600 29.200 ;
        RECT 139.000 26.800 139.400 27.200 ;
        RECT 140.600 25.800 141.000 26.200 ;
        RECT 136.600 24.800 137.000 25.200 ;
        RECT 136.600 24.200 136.900 24.800 ;
        RECT 136.600 23.800 137.000 24.200 ;
        RECT 137.400 22.800 137.800 23.200 ;
        RECT 136.600 21.800 137.000 22.200 ;
        RECT 136.600 19.200 136.900 21.800 ;
        RECT 136.600 18.800 137.000 19.200 ;
        RECT 127.000 13.800 127.400 14.200 ;
        RECT 119.000 12.800 120.200 13.100 ;
        RECT 107.000 11.800 108.100 12.100 ;
        RECT 112.600 11.800 113.000 12.200 ;
        RECT 96.600 9.800 97.000 10.200 ;
        RECT 96.600 9.200 96.900 9.800 ;
        RECT 107.000 9.200 107.300 11.800 ;
        RECT 83.800 8.800 84.200 9.200 ;
        RECT 95.000 8.800 95.400 9.200 ;
        RECT 96.600 8.800 97.000 9.200 ;
        RECT 83.000 6.800 83.400 7.200 ;
        RECT 86.200 6.800 86.600 7.200 ;
        RECT 90.200 6.800 90.600 7.200 ;
        RECT 86.200 6.200 86.500 6.800 ;
        RECT 90.200 6.200 90.500 6.800 ;
        RECT 86.200 5.800 86.600 6.200 ;
        RECT 89.400 5.800 89.800 6.200 ;
        RECT 90.200 5.800 90.600 6.200 ;
        RECT 92.600 6.100 93.000 6.200 ;
        RECT 93.400 6.100 93.800 6.200 ;
        RECT 92.600 5.800 93.800 6.100 ;
        RECT 89.400 5.200 89.700 5.800 ;
        RECT 89.400 4.800 89.800 5.200 ;
        RECT 99.000 3.100 99.400 8.900 ;
        RECT 102.200 6.200 102.600 6.300 ;
        RECT 103.000 6.200 103.400 6.300 ;
        RECT 102.200 5.900 103.400 6.200 ;
        RECT 103.800 3.100 104.200 8.900 ;
        RECT 104.600 8.800 105.000 9.200 ;
        RECT 107.000 8.800 107.400 9.200 ;
        RECT 104.600 7.200 104.900 8.800 ;
        RECT 104.600 6.800 105.000 7.200 ;
        RECT 105.400 5.100 105.800 7.900 ;
        RECT 108.600 5.100 109.000 7.900 ;
        RECT 110.200 3.100 110.600 8.900 ;
        RECT 111.800 8.800 112.200 9.200 ;
        RECT 111.800 7.200 112.100 8.800 ;
        RECT 111.800 6.800 112.200 7.200 ;
        RECT 112.600 6.200 112.900 11.800 ;
        RECT 113.400 10.200 113.700 12.800 ;
        RECT 116.600 11.800 117.000 12.200 ;
        RECT 113.400 9.800 113.800 10.200 ;
        RECT 112.600 5.800 113.000 6.200 ;
        RECT 115.000 3.100 115.400 8.900 ;
        RECT 116.600 6.200 116.900 11.800 ;
        RECT 117.400 9.200 117.700 12.800 ;
        RECT 123.000 12.100 123.400 12.200 ;
        RECT 123.800 12.100 124.200 12.200 ;
        RECT 123.000 11.800 124.200 12.100 ;
        RECT 123.000 10.800 123.400 11.200 ;
        RECT 123.000 9.200 123.300 10.800 ;
        RECT 127.000 9.200 127.300 13.800 ;
        RECT 127.800 12.100 128.200 17.900 ;
        RECT 129.400 15.100 129.800 15.200 ;
        RECT 130.200 15.100 130.600 15.200 ;
        RECT 129.400 14.800 130.600 15.100 ;
        RECT 132.600 12.100 133.000 17.900 ;
        RECT 136.600 16.800 137.000 17.200 ;
        RECT 136.600 9.200 136.900 16.800 ;
        RECT 117.400 8.800 117.800 9.200 ;
        RECT 123.000 8.800 123.400 9.200 ;
        RECT 127.000 8.800 127.400 9.200 ;
        RECT 116.600 5.800 117.000 6.200 ;
        RECT 121.400 6.100 121.800 6.200 ;
        RECT 122.200 6.100 122.600 6.200 ;
        RECT 121.400 5.800 122.600 6.100 ;
        RECT 126.200 5.100 126.600 7.900 ;
        RECT 127.000 7.200 127.300 8.800 ;
        RECT 127.000 6.800 127.400 7.200 ;
        RECT 127.800 3.100 128.200 8.900 ;
        RECT 129.400 7.800 129.800 8.200 ;
        RECT 129.400 6.200 129.700 7.800 ;
        RECT 129.400 5.800 129.800 6.200 ;
        RECT 132.600 3.100 133.000 8.900 ;
        RECT 136.600 8.800 137.000 9.200 ;
        RECT 135.800 7.800 136.200 8.200 ;
        RECT 135.800 7.200 136.100 7.800 ;
        RECT 135.800 6.800 136.200 7.200 ;
        RECT 137.400 5.200 137.700 22.800 ;
        RECT 140.600 18.200 140.900 25.800 ;
        RECT 141.400 24.800 141.800 25.200 ;
        RECT 141.400 23.200 141.700 24.800 ;
        RECT 141.400 22.800 141.800 23.200 ;
        RECT 140.600 17.800 141.000 18.200 ;
        RECT 140.600 16.800 141.000 17.200 ;
        RECT 140.600 15.200 140.900 16.800 ;
        RECT 143.000 15.200 143.300 30.800 ;
        RECT 143.800 28.800 144.200 29.200 ;
        RECT 144.600 29.100 145.000 29.200 ;
        RECT 145.400 29.100 145.800 29.200 ;
        RECT 144.600 28.800 145.800 29.100 ;
        RECT 143.800 28.200 144.100 28.800 ;
        RECT 143.800 27.800 144.200 28.200 ;
        RECT 146.200 28.100 146.500 34.800 ;
        RECT 147.000 33.800 147.400 34.200 ;
        RECT 147.000 32.200 147.300 33.800 ;
        RECT 147.800 33.100 148.200 35.900 ;
        RECT 147.000 31.800 147.400 32.200 ;
        RECT 145.400 27.800 146.500 28.100 ;
        RECT 145.400 22.200 145.700 27.800 ;
        RECT 146.200 24.800 146.600 25.200 ;
        RECT 144.600 21.800 145.000 22.200 ;
        RECT 145.400 21.800 145.800 22.200 ;
        RECT 144.600 15.200 144.900 21.800 ;
        RECT 146.200 19.200 146.500 24.800 ;
        RECT 147.800 23.100 148.200 28.900 ;
        RECT 146.200 18.800 146.600 19.200 ;
        RECT 148.600 17.200 148.900 38.800 ;
        RECT 149.400 32.100 149.800 37.900 ;
        RECT 150.200 34.200 150.500 45.800 ;
        RECT 151.000 41.800 151.400 42.200 ;
        RECT 151.000 35.200 151.300 41.800 ;
        RECT 151.800 40.200 152.100 45.800 ;
        RECT 151.800 39.800 152.200 40.200 ;
        RECT 151.000 34.800 151.400 35.200 ;
        RECT 150.200 33.800 150.600 34.200 ;
        RECT 153.400 32.200 153.700 46.800 ;
        RECT 154.200 45.800 154.600 46.200 ;
        RECT 154.200 45.200 154.500 45.800 ;
        RECT 154.200 44.800 154.600 45.200 ;
        RECT 153.400 31.800 153.800 32.200 ;
        RECT 154.200 32.100 154.600 37.900 ;
        RECT 149.400 26.100 149.800 26.200 ;
        RECT 150.200 26.100 150.600 26.200 ;
        RECT 149.400 25.800 150.600 26.100 ;
        RECT 151.000 25.800 151.400 26.200 ;
        RECT 151.000 25.200 151.300 25.800 ;
        RECT 151.000 24.800 151.400 25.200 ;
        RECT 152.600 23.100 153.000 28.900 ;
        RECT 153.400 27.200 153.700 31.800 ;
        RECT 155.000 28.200 155.300 50.800 ;
        RECT 155.800 49.200 156.100 53.800 ;
        RECT 156.600 51.800 157.000 52.200 ;
        RECT 156.600 51.200 156.900 51.800 ;
        RECT 156.600 50.800 157.000 51.200 ;
        RECT 156.600 49.800 157.000 50.200 ;
        RECT 156.600 49.200 156.900 49.800 ;
        RECT 155.800 48.800 156.200 49.200 ;
        RECT 156.600 48.800 157.000 49.200 ;
        RECT 155.800 45.100 156.200 45.200 ;
        RECT 155.800 44.800 156.900 45.100 ;
        RECT 155.800 43.800 156.200 44.200 ;
        RECT 155.800 29.200 156.100 43.800 ;
        RECT 156.600 29.200 156.900 44.800 ;
        RECT 158.200 44.200 158.500 65.800 ;
        RECT 159.800 64.200 160.100 85.800 ;
        RECT 162.200 85.800 162.600 86.200 ;
        RECT 165.400 86.100 165.800 86.200 ;
        RECT 164.600 85.800 165.800 86.100 ;
        RECT 167.000 85.800 167.400 86.200 ;
        RECT 162.200 85.200 162.500 85.800 ;
        RECT 162.200 84.800 162.600 85.200 ;
        RECT 162.200 74.800 162.600 75.200 ;
        RECT 162.200 66.200 162.500 74.800 ;
        RECT 163.800 71.800 164.200 72.200 ;
        RECT 163.800 71.200 164.100 71.800 ;
        RECT 163.800 70.800 164.200 71.200 ;
        RECT 163.800 68.800 164.200 69.200 ;
        RECT 163.000 67.800 163.400 68.200 ;
        RECT 163.000 67.200 163.300 67.800 ;
        RECT 163.000 66.800 163.400 67.200 ;
        RECT 163.800 66.200 164.100 68.800 ;
        RECT 164.600 66.200 164.900 85.800 ;
        RECT 167.000 84.200 167.300 85.800 ;
        RECT 167.000 83.800 167.400 84.200 ;
        RECT 165.400 75.800 165.800 76.200 ;
        RECT 165.400 75.200 165.700 75.800 ;
        RECT 165.400 74.800 165.800 75.200 ;
        RECT 166.200 74.800 166.600 75.200 ;
        RECT 166.200 74.200 166.500 74.800 ;
        RECT 166.200 73.800 166.600 74.200 ;
        RECT 167.000 68.800 167.400 69.200 ;
        RECT 167.000 68.200 167.300 68.800 ;
        RECT 167.000 67.800 167.400 68.200 ;
        RECT 167.800 67.200 168.100 86.800 ;
        RECT 168.600 86.200 168.900 86.800 ;
        RECT 171.000 86.200 171.300 87.800 ;
        RECT 168.600 85.800 169.000 86.200 ;
        RECT 169.400 86.100 169.800 86.200 ;
        RECT 170.200 86.100 170.600 86.200 ;
        RECT 169.400 85.800 170.600 86.100 ;
        RECT 171.000 85.800 171.400 86.200 ;
        RECT 169.400 75.200 169.700 85.800 ;
        RECT 171.800 85.200 172.100 115.800 ;
        RECT 173.400 114.800 173.800 115.200 ;
        RECT 173.400 113.200 173.700 114.800 ;
        RECT 173.400 112.800 173.800 113.200 ;
        RECT 174.200 112.800 174.600 113.200 ;
        RECT 174.200 111.200 174.500 112.800 ;
        RECT 175.000 112.200 175.300 121.800 ;
        RECT 175.000 111.800 175.400 112.200 ;
        RECT 174.200 110.800 174.600 111.200 ;
        RECT 172.600 103.800 173.000 104.200 ;
        RECT 172.600 99.100 172.900 103.800 ;
        RECT 173.400 103.100 173.800 108.900 ;
        RECT 176.600 107.200 176.900 125.800 ;
        RECT 177.400 123.100 177.800 128.900 ;
        RECT 179.800 124.200 180.100 132.800 ;
        RECT 179.800 123.800 180.200 124.200 ;
        RECT 179.800 121.800 180.200 122.200 ;
        RECT 179.800 121.200 180.100 121.800 ;
        RECT 179.800 120.800 180.200 121.200 ;
        RECT 176.600 106.800 177.000 107.200 ;
        RECT 175.800 106.100 176.200 106.200 ;
        RECT 176.600 106.100 177.000 106.200 ;
        RECT 175.800 105.800 177.000 106.100 ;
        RECT 178.200 103.100 178.600 108.900 ;
        RECT 179.800 105.100 180.200 107.900 ;
        RECT 172.600 98.800 173.700 99.100 ;
        RECT 172.600 92.100 173.000 97.900 ;
        RECT 173.400 94.200 173.700 98.800 ;
        RECT 173.400 93.800 173.800 94.200 ;
        RECT 174.200 93.100 174.600 95.900 ;
        RECT 175.000 94.800 175.400 95.200 ;
        RECT 177.400 94.800 177.800 95.200 ;
        RECT 175.000 93.200 175.300 94.800 ;
        RECT 175.000 92.800 175.400 93.200 ;
        RECT 173.400 91.800 173.800 92.200 ;
        RECT 173.400 89.200 173.700 91.800 ;
        RECT 177.400 91.200 177.700 94.800 ;
        RECT 177.400 90.800 177.800 91.200 ;
        RECT 173.400 88.800 173.800 89.200 ;
        RECT 172.600 88.100 173.000 88.200 ;
        RECT 173.400 88.100 173.800 88.200 ;
        RECT 172.600 87.800 173.800 88.100 ;
        RECT 179.800 87.800 180.200 88.200 ;
        RECT 178.200 86.800 178.600 87.200 ;
        RECT 178.200 86.200 178.500 86.800 ;
        RECT 178.200 85.800 178.600 86.200 ;
        RECT 170.200 85.100 170.600 85.200 ;
        RECT 171.000 85.100 171.400 85.200 ;
        RECT 170.200 84.800 171.400 85.100 ;
        RECT 171.800 84.800 172.200 85.200 ;
        RECT 170.200 79.100 170.600 79.200 ;
        RECT 171.000 79.100 171.400 79.200 ;
        RECT 170.200 78.800 171.400 79.100 ;
        RECT 168.600 74.800 169.000 75.200 ;
        RECT 169.400 74.800 169.800 75.200 ;
        RECT 168.600 74.200 168.900 74.800 ;
        RECT 168.600 73.800 169.000 74.200 ;
        RECT 168.600 71.800 169.000 72.200 ;
        RECT 172.600 72.100 173.000 77.900 ;
        RECT 175.000 75.100 175.400 75.200 ;
        RECT 175.800 75.100 176.200 75.200 ;
        RECT 175.000 74.800 176.200 75.100 ;
        RECT 175.800 73.800 176.200 74.200 ;
        RECT 168.600 68.200 168.900 71.800 ;
        RECT 168.600 67.800 169.000 68.200 ;
        RECT 166.200 66.800 166.600 67.200 ;
        RECT 167.800 66.800 168.200 67.200 ;
        RECT 160.600 66.100 161.000 66.200 ;
        RECT 161.400 66.100 161.800 66.200 ;
        RECT 160.600 65.800 161.800 66.100 ;
        RECT 162.200 65.800 162.600 66.200 ;
        RECT 163.800 65.800 164.200 66.200 ;
        RECT 164.600 66.100 165.000 66.200 ;
        RECT 165.400 66.100 165.800 66.200 ;
        RECT 164.600 65.800 165.800 66.100 ;
        RECT 159.800 63.800 160.200 64.200 ;
        RECT 159.800 61.800 160.200 62.200 ;
        RECT 159.800 58.200 160.100 61.800 ;
        RECT 161.400 59.800 161.800 60.200 ;
        RECT 159.800 57.800 160.200 58.200 ;
        RECT 161.400 55.200 161.700 59.800 ;
        RECT 161.400 54.800 161.800 55.200 ;
        RECT 160.600 54.100 161.000 54.200 ;
        RECT 161.400 54.100 161.800 54.200 ;
        RECT 160.600 53.800 161.800 54.100 ;
        RECT 159.800 52.800 160.200 53.200 ;
        RECT 158.200 43.800 158.600 44.200 ;
        RECT 159.000 43.100 159.400 48.900 ;
        RECT 159.800 48.200 160.100 52.800 ;
        RECT 161.400 50.800 161.800 51.200 ;
        RECT 159.800 47.800 160.200 48.200 ;
        RECT 159.800 46.800 160.200 47.200 ;
        RECT 159.800 46.200 160.100 46.800 ;
        RECT 161.400 46.200 161.700 50.800 ;
        RECT 159.800 45.800 160.200 46.200 ;
        RECT 161.400 45.800 161.800 46.200 ;
        RECT 162.200 42.200 162.500 65.800 ;
        RECT 163.000 63.800 163.400 64.200 ;
        RECT 163.000 56.100 163.300 63.800 ;
        RECT 163.800 61.800 164.200 62.200 ;
        RECT 163.800 60.200 164.100 61.800 ;
        RECT 163.800 59.800 164.200 60.200 ;
        RECT 163.000 55.700 163.400 56.100 ;
        RECT 165.400 55.800 165.800 56.200 ;
        RECT 165.400 55.200 165.700 55.800 ;
        RECT 166.200 55.200 166.500 66.800 ;
        RECT 167.000 65.800 167.400 66.200 ;
        RECT 167.800 65.800 168.200 66.200 ;
        RECT 167.000 65.200 167.300 65.800 ;
        RECT 167.000 64.800 167.400 65.200 ;
        RECT 167.800 59.200 168.100 65.800 ;
        RECT 171.800 63.100 172.200 68.900 ;
        RECT 175.800 68.200 176.100 73.800 ;
        RECT 177.400 72.100 177.800 77.900 ;
        RECT 179.000 73.100 179.400 75.900 ;
        RECT 179.800 69.200 180.100 87.800 ;
        RECT 175.800 67.800 176.200 68.200 ;
        RECT 174.200 66.800 174.600 67.200 ;
        RECT 172.600 66.100 173.000 66.200 ;
        RECT 173.400 66.100 173.800 66.200 ;
        RECT 172.600 65.800 173.800 66.100 ;
        RECT 169.400 62.100 169.800 62.200 ;
        RECT 170.200 62.100 170.600 62.200 ;
        RECT 169.400 61.800 170.600 62.100 ;
        RECT 169.400 60.800 169.800 61.200 ;
        RECT 167.800 58.800 168.200 59.200 ;
        RECT 168.600 56.800 169.000 57.200 ;
        RECT 168.600 55.200 168.900 56.800 ;
        RECT 165.400 54.800 165.800 55.200 ;
        RECT 166.200 54.800 166.600 55.200 ;
        RECT 168.600 54.800 169.000 55.200 ;
        RECT 166.200 49.200 166.500 54.800 ;
        RECT 168.600 53.800 169.000 54.200 ;
        RECT 168.600 49.200 168.900 53.800 ;
        RECT 169.400 49.200 169.700 60.800 ;
        RECT 170.200 59.100 170.600 59.200 ;
        RECT 171.000 59.100 171.400 59.200 ;
        RECT 170.200 58.800 171.400 59.100 ;
        RECT 170.200 55.800 170.600 56.200 ;
        RECT 163.800 43.100 164.200 48.900 ;
        RECT 166.200 48.800 166.600 49.200 ;
        RECT 168.600 48.800 169.000 49.200 ;
        RECT 169.400 48.800 169.800 49.200 ;
        RECT 170.200 48.200 170.500 55.800 ;
        RECT 172.600 52.100 173.000 57.900 ;
        RECT 174.200 55.200 174.500 66.800 ;
        RECT 176.600 63.100 177.000 68.900 ;
        RECT 179.800 68.800 180.200 69.200 ;
        RECT 178.200 65.100 178.600 67.900 ;
        RECT 179.000 67.800 179.400 68.200 ;
        RECT 179.000 58.200 179.300 67.800 ;
        RECT 179.800 61.800 180.200 62.200 ;
        RECT 174.200 54.800 174.600 55.200 ;
        RECT 165.400 45.100 165.800 47.900 ;
        RECT 166.200 47.800 166.600 48.200 ;
        RECT 170.200 47.800 170.600 48.200 ;
        RECT 166.200 47.200 166.500 47.800 ;
        RECT 166.200 46.800 166.600 47.200 ;
        RECT 168.600 46.800 169.000 47.200 ;
        RECT 167.000 45.800 167.400 46.200 ;
        RECT 162.200 41.800 162.600 42.200 ;
        RECT 163.000 40.800 163.400 41.200 ;
        RECT 164.600 40.800 165.000 41.200 ;
        RECT 158.200 39.800 158.600 40.200 ;
        RECT 158.200 39.200 158.500 39.800 ;
        RECT 158.200 38.800 158.600 39.200 ;
        RECT 161.400 35.100 161.800 35.200 ;
        RECT 162.200 35.100 162.600 35.200 ;
        RECT 161.400 34.800 162.600 35.100 ;
        RECT 159.000 33.100 159.400 33.200 ;
        RECT 158.200 32.800 159.400 33.100 ;
        RECT 155.800 28.800 156.200 29.200 ;
        RECT 156.600 28.800 157.000 29.200 ;
        RECT 153.400 26.800 153.800 27.200 ;
        RECT 154.200 25.100 154.600 27.900 ;
        RECT 155.000 27.800 155.400 28.200 ;
        RECT 158.200 27.200 158.500 32.800 ;
        RECT 159.000 32.200 159.300 32.800 ;
        RECT 159.000 31.800 159.400 32.200 ;
        RECT 159.800 27.800 160.200 28.200 ;
        RECT 158.200 26.800 158.600 27.200 ;
        RECT 158.200 25.800 158.600 26.200 ;
        RECT 156.600 24.800 157.000 25.200 ;
        RECT 156.600 23.200 156.900 24.800 ;
        RECT 156.600 22.800 157.000 23.200 ;
        RECT 152.600 17.800 153.000 18.200 ;
        RECT 147.000 16.800 147.400 17.200 ;
        RECT 148.600 16.800 149.000 17.200 ;
        RECT 147.000 15.200 147.300 16.800 ;
        RECT 148.600 15.800 149.000 16.200 ;
        RECT 148.600 15.200 148.900 15.800 ;
        RECT 152.600 15.200 152.900 17.800 ;
        RECT 138.200 14.800 138.600 15.200 ;
        RECT 140.600 14.800 141.000 15.200 ;
        RECT 143.000 14.800 143.400 15.200 ;
        RECT 144.600 14.800 145.000 15.200 ;
        RECT 147.000 14.800 147.400 15.200 ;
        RECT 147.800 14.800 148.200 15.200 ;
        RECT 148.600 14.800 149.000 15.200 ;
        RECT 149.400 14.800 149.800 15.200 ;
        RECT 151.800 14.800 152.200 15.200 ;
        RECT 152.600 14.800 153.000 15.200 ;
        RECT 138.200 14.200 138.500 14.800 ;
        RECT 147.800 14.200 148.100 14.800 ;
        RECT 138.200 13.800 138.600 14.200 ;
        RECT 146.200 13.800 146.600 14.200 ;
        RECT 147.800 13.800 148.200 14.200 ;
        RECT 144.600 12.800 145.000 13.200 ;
        RECT 138.200 8.800 138.600 9.200 ;
        RECT 138.200 8.200 138.500 8.800 ;
        RECT 138.200 7.800 138.600 8.200 ;
        RECT 140.600 8.100 141.000 8.200 ;
        RECT 139.800 7.800 141.000 8.100 ;
        RECT 139.800 7.200 140.100 7.800 ;
        RECT 139.800 6.800 140.200 7.200 ;
        RECT 144.600 6.200 144.900 12.800 ;
        RECT 146.200 7.200 146.500 13.800 ;
        RECT 149.400 13.200 149.700 14.800 ;
        RECT 151.800 14.200 152.100 14.800 ;
        RECT 151.800 13.800 152.200 14.200 ;
        RECT 149.400 12.800 149.800 13.200 ;
        RECT 153.400 13.100 153.800 15.900 ;
        RECT 154.200 13.800 154.600 14.200 ;
        RECT 146.200 6.800 146.600 7.200 ;
        RECT 149.400 7.100 149.800 7.200 ;
        RECT 150.200 7.100 150.600 7.200 ;
        RECT 149.400 6.800 150.600 7.100 ;
        RECT 146.200 6.200 146.500 6.800 ;
        RECT 143.800 6.100 144.200 6.200 ;
        RECT 144.600 6.100 145.000 6.200 ;
        RECT 143.800 5.800 145.000 6.100 ;
        RECT 146.200 5.800 146.600 6.200 ;
        RECT 147.000 5.800 147.400 6.200 ;
        RECT 149.400 6.100 149.800 6.200 ;
        RECT 150.200 6.100 150.600 6.200 ;
        RECT 149.400 5.800 150.600 6.100 ;
        RECT 147.000 5.200 147.300 5.800 ;
        RECT 137.400 4.800 137.800 5.200 ;
        RECT 147.000 4.800 147.400 5.200 ;
        RECT 151.000 5.100 151.400 7.900 ;
        RECT 152.600 3.100 153.000 8.900 ;
        RECT 154.200 7.200 154.500 13.800 ;
        RECT 155.000 12.100 155.400 17.900 ;
        RECT 155.800 15.800 156.200 16.200 ;
        RECT 155.800 15.100 156.100 15.800 ;
        RECT 158.200 15.200 158.500 25.800 ;
        RECT 159.000 21.800 159.400 22.200 ;
        RECT 159.000 18.200 159.300 21.800 ;
        RECT 159.800 19.200 160.100 27.800 ;
        RECT 160.600 25.100 161.000 27.900 ;
        RECT 161.400 26.800 161.800 27.200 ;
        RECT 161.400 26.200 161.700 26.800 ;
        RECT 161.400 25.800 161.800 26.200 ;
        RECT 159.800 18.800 160.200 19.200 ;
        RECT 159.000 17.800 159.400 18.200 ;
        RECT 155.800 14.700 156.200 15.100 ;
        RECT 158.200 14.800 158.600 15.200 ;
        RECT 159.800 12.100 160.200 17.900 ;
        RECT 159.800 9.100 160.200 9.200 ;
        RECT 160.600 9.100 161.000 9.200 ;
        RECT 153.400 6.800 153.800 7.200 ;
        RECT 154.200 6.800 154.600 7.200 ;
        RECT 153.400 6.300 153.700 6.800 ;
        RECT 153.400 5.900 153.800 6.300 ;
        RECT 157.400 3.100 157.800 8.900 ;
        RECT 159.800 8.800 161.000 9.100 ;
        RECT 160.600 5.100 161.000 7.900 ;
        RECT 161.400 7.200 161.700 25.800 ;
        RECT 162.200 23.100 162.600 28.900 ;
        RECT 162.200 19.800 162.600 20.200 ;
        RECT 162.200 19.200 162.500 19.800 ;
        RECT 162.200 18.800 162.600 19.200 ;
        RECT 163.000 15.200 163.300 40.800 ;
        RECT 163.800 35.800 164.200 36.200 ;
        RECT 163.800 35.200 164.100 35.800 ;
        RECT 164.600 35.200 164.900 40.800 ;
        RECT 167.000 40.200 167.300 45.800 ;
        RECT 168.600 45.200 168.900 46.800 ;
        RECT 169.400 45.800 169.800 46.200 ;
        RECT 169.400 45.200 169.700 45.800 ;
        RECT 168.600 44.800 169.000 45.200 ;
        RECT 169.400 44.800 169.800 45.200 ;
        RECT 167.000 39.800 167.400 40.200 ;
        RECT 163.800 34.800 164.200 35.200 ;
        RECT 164.600 34.800 165.000 35.200 ;
        RECT 164.600 32.100 165.000 32.200 ;
        RECT 165.400 32.100 165.800 32.200 ;
        RECT 167.800 32.100 168.200 37.900 ;
        RECT 169.400 35.200 169.700 44.800 ;
        RECT 173.400 43.100 173.800 48.900 ;
        RECT 174.200 46.200 174.500 54.800 ;
        RECT 176.600 54.700 177.000 55.100 ;
        RECT 176.600 54.200 176.900 54.700 ;
        RECT 176.600 53.800 177.000 54.200 ;
        RECT 175.000 51.800 175.400 52.200 ;
        RECT 177.400 52.100 177.800 57.900 ;
        RECT 179.000 57.800 179.400 58.200 ;
        RECT 179.000 53.100 179.400 55.900 ;
        RECT 174.200 45.800 174.600 46.200 ;
        RECT 174.200 45.200 174.500 45.800 ;
        RECT 174.200 44.800 174.600 45.200 ;
        RECT 171.000 42.100 171.400 42.200 ;
        RECT 171.800 42.100 172.200 42.200 ;
        RECT 171.000 41.800 172.200 42.100 ;
        RECT 171.800 39.800 172.200 40.200 ;
        RECT 169.400 34.800 169.800 35.200 ;
        RECT 170.200 35.100 170.600 35.200 ;
        RECT 171.000 35.100 171.400 35.200 ;
        RECT 170.200 34.800 171.400 35.100 ;
        RECT 164.600 31.800 165.800 32.100 ;
        RECT 169.400 30.200 169.700 34.800 ;
        RECT 170.200 33.800 170.600 34.200 ;
        RECT 169.400 29.800 169.800 30.200 ;
        RECT 170.200 29.200 170.500 33.800 ;
        RECT 171.000 32.800 171.400 33.200 ;
        RECT 164.600 25.800 165.000 26.200 ;
        RECT 164.600 19.200 164.900 25.800 ;
        RECT 167.000 23.100 167.400 28.900 ;
        RECT 169.400 28.800 169.800 29.200 ;
        RECT 170.200 28.800 170.600 29.200 ;
        RECT 169.400 28.200 169.700 28.800 ;
        RECT 171.000 28.200 171.300 32.800 ;
        RECT 171.800 29.200 172.100 39.800 ;
        RECT 172.600 32.100 173.000 37.900 ;
        RECT 174.200 33.100 174.600 35.900 ;
        RECT 175.000 35.200 175.300 51.800 ;
        RECT 177.400 50.800 177.800 51.200 ;
        RECT 175.800 46.100 176.200 46.200 ;
        RECT 176.600 46.100 177.000 46.200 ;
        RECT 175.800 45.800 177.000 46.100 ;
        RECT 176.600 43.800 177.000 44.200 ;
        RECT 176.600 39.200 176.900 43.800 ;
        RECT 176.600 38.800 177.000 39.200 ;
        RECT 175.800 35.800 176.200 36.200 ;
        RECT 175.800 35.200 176.100 35.800 ;
        RECT 175.000 34.800 175.400 35.200 ;
        RECT 175.800 34.800 176.200 35.200 ;
        RECT 177.400 29.200 177.700 50.800 ;
        RECT 179.800 49.100 180.100 61.800 ;
        RECT 178.200 43.100 178.600 48.900 ;
        RECT 179.000 48.800 180.100 49.100 ;
        RECT 178.200 36.800 178.600 37.200 ;
        RECT 178.200 35.200 178.500 36.800 ;
        RECT 178.200 34.800 178.600 35.200 ;
        RECT 171.800 28.800 172.200 29.200 ;
        RECT 177.400 28.800 177.800 29.200 ;
        RECT 169.400 27.800 169.800 28.200 ;
        RECT 171.000 27.800 171.400 28.200 ;
        RECT 173.400 27.100 173.800 27.200 ;
        RECT 174.200 27.100 174.600 27.200 ;
        RECT 173.400 26.800 174.600 27.100 ;
        RECT 179.000 26.200 179.300 48.800 ;
        RECT 179.800 45.100 180.200 47.900 ;
        RECT 179.800 28.800 180.200 29.200 ;
        RECT 179.800 27.200 180.100 28.800 ;
        RECT 179.800 26.800 180.200 27.200 ;
        RECT 173.400 26.100 173.800 26.200 ;
        RECT 174.200 26.100 174.600 26.200 ;
        RECT 173.400 25.800 174.600 26.100 ;
        RECT 175.800 25.800 176.200 26.200 ;
        RECT 179.000 25.800 179.400 26.200 ;
        RECT 171.800 24.800 172.200 25.200 ;
        RECT 173.400 24.800 173.800 25.200 ;
        RECT 171.800 24.200 172.100 24.800 ;
        RECT 168.600 23.800 169.000 24.200 ;
        RECT 171.800 23.800 172.200 24.200 ;
        RECT 168.600 19.200 168.900 23.800 ;
        RECT 169.400 22.800 169.800 23.200 ;
        RECT 169.400 22.200 169.700 22.800 ;
        RECT 169.400 21.800 169.800 22.200 ;
        RECT 164.600 18.800 165.000 19.200 ;
        RECT 168.600 18.800 169.000 19.200 ;
        RECT 169.400 16.200 169.700 21.800 ;
        RECT 173.400 19.200 173.700 24.800 ;
        RECT 174.200 22.800 174.600 23.200 ;
        RECT 173.400 18.800 173.800 19.200 ;
        RECT 166.200 15.800 166.600 16.200 ;
        RECT 169.400 15.800 169.800 16.200 ;
        RECT 170.200 16.100 170.600 16.200 ;
        RECT 171.000 16.100 171.400 16.200 ;
        RECT 170.200 15.800 171.400 16.100 ;
        RECT 171.800 16.100 172.200 16.200 ;
        RECT 172.600 16.100 173.000 16.200 ;
        RECT 171.800 15.800 173.000 16.100 ;
        RECT 166.200 15.200 166.500 15.800 ;
        RECT 163.000 14.800 163.400 15.200 ;
        RECT 163.800 15.100 164.200 15.200 ;
        RECT 164.600 15.100 165.000 15.200 ;
        RECT 163.800 14.800 165.000 15.100 ;
        RECT 166.200 14.800 166.600 15.200 ;
        RECT 163.000 14.200 163.300 14.800 ;
        RECT 163.000 13.800 163.400 14.200 ;
        RECT 167.800 13.800 168.200 14.200 ;
        RECT 163.800 10.800 164.200 11.200 ;
        RECT 161.400 6.800 161.800 7.200 ;
        RECT 162.200 3.100 162.600 8.900 ;
        RECT 163.800 6.200 164.100 10.800 ;
        RECT 167.800 9.200 168.100 13.800 ;
        RECT 174.200 13.200 174.500 22.800 ;
        RECT 175.800 16.200 176.100 25.800 ;
        RECT 178.200 24.800 178.600 25.200 ;
        RECT 178.200 22.200 178.500 24.800 ;
        RECT 178.200 21.800 178.600 22.200 ;
        RECT 179.000 16.800 179.400 17.200 ;
        RECT 175.800 15.800 176.200 16.200 ;
        RECT 175.800 15.200 176.100 15.800 ;
        RECT 179.000 15.200 179.300 16.800 ;
        RECT 175.800 14.800 176.200 15.200 ;
        RECT 177.400 15.100 177.800 15.200 ;
        RECT 178.200 15.100 178.600 15.200 ;
        RECT 177.400 14.800 178.600 15.100 ;
        RECT 179.000 14.800 179.400 15.200 ;
        RECT 170.200 13.100 170.600 13.200 ;
        RECT 171.000 13.100 171.400 13.200 ;
        RECT 170.200 12.800 171.400 13.100 ;
        RECT 171.800 12.800 172.200 13.200 ;
        RECT 174.200 12.800 174.600 13.200 ;
        RECT 171.800 10.200 172.100 12.800 ;
        RECT 176.600 11.800 177.000 12.200 ;
        RECT 176.600 11.200 176.900 11.800 ;
        RECT 176.600 10.800 177.000 11.200 ;
        RECT 169.400 9.800 169.800 10.200 ;
        RECT 171.800 9.800 172.200 10.200 ;
        RECT 179.000 9.800 179.400 10.200 ;
        RECT 169.400 9.200 169.700 9.800 ;
        RECT 179.000 9.200 179.300 9.800 ;
        RECT 163.800 5.800 164.200 6.200 ;
        RECT 167.000 3.100 167.400 8.900 ;
        RECT 167.800 8.800 168.200 9.200 ;
        RECT 169.400 8.800 169.800 9.200 ;
        RECT 170.200 5.100 170.600 7.900 ;
        RECT 171.000 7.800 171.400 8.200 ;
        RECT 171.000 7.200 171.300 7.800 ;
        RECT 171.000 6.800 171.400 7.200 ;
        RECT 171.800 3.100 172.200 8.900 ;
        RECT 172.600 6.800 173.000 7.200 ;
        RECT 172.600 6.300 172.900 6.800 ;
        RECT 172.600 5.900 173.000 6.300 ;
        RECT 176.600 3.100 177.000 8.900 ;
        RECT 179.000 8.800 179.400 9.200 ;
      LAYER via2 ;
        RECT 19.000 155.800 19.400 156.200 ;
        RECT 20.600 154.800 21.000 155.200 ;
        RECT 12.600 153.800 13.000 154.200 ;
        RECT 11.000 152.800 11.400 153.200 ;
        RECT 4.600 145.800 5.000 146.200 ;
        RECT 11.000 147.800 11.400 148.200 ;
        RECT 14.200 134.800 14.600 135.200 ;
        RECT 2.200 125.800 2.600 126.200 ;
        RECT 2.200 114.800 2.600 115.200 ;
        RECT 2.200 54.800 2.600 55.200 ;
        RECT 19.800 136.800 20.200 137.200 ;
        RECT 23.000 134.800 23.400 135.200 ;
        RECT 54.200 165.800 54.600 166.200 ;
        RECT 54.200 157.800 54.600 158.200 ;
        RECT 40.600 146.800 41.000 147.200 ;
        RECT 42.200 144.800 42.600 145.200 ;
        RECT 34.200 136.800 34.600 137.200 ;
        RECT 27.800 134.800 28.200 135.200 ;
        RECT 33.400 134.800 33.800 135.200 ;
        RECT 39.000 132.800 39.400 133.200 ;
        RECT 18.200 113.800 18.600 114.200 ;
        RECT 11.800 106.800 12.200 107.200 ;
        RECT 12.600 105.800 13.000 106.200 ;
        RECT 25.400 123.800 25.800 124.200 ;
        RECT 35.800 128.800 36.200 129.200 ;
        RECT 10.200 88.800 10.600 89.200 ;
        RECT 11.000 87.800 11.400 88.200 ;
        RECT 21.400 94.800 21.800 95.200 ;
        RECT 14.200 87.800 14.600 88.200 ;
        RECT 18.200 84.800 18.600 85.200 ;
        RECT 10.200 68.800 10.600 69.200 ;
        RECT 15.000 72.800 15.400 73.200 ;
        RECT 22.200 86.800 22.600 87.200 ;
        RECT 39.000 125.800 39.400 126.200 ;
        RECT 34.200 112.800 34.600 113.200 ;
        RECT 26.200 85.800 26.600 86.200 ;
        RECT 27.800 84.800 28.200 85.200 ;
        RECT 30.200 74.800 30.600 75.200 ;
        RECT 39.000 108.800 39.400 109.200 ;
        RECT 38.200 96.800 38.600 97.200 ;
        RECT 50.200 151.800 50.600 152.200 ;
        RECT 60.600 155.800 61.000 156.200 ;
        RECT 102.200 165.800 102.600 166.200 ;
        RECT 56.600 148.800 57.000 149.200 ;
        RECT 50.200 134.800 50.600 135.200 ;
        RECT 49.400 131.800 49.800 132.200 ;
        RECT 83.000 154.700 83.400 155.100 ;
        RECT 93.400 158.800 93.800 159.200 ;
        RECT 82.200 145.800 82.600 146.200 ;
        RECT 66.200 125.800 66.600 126.200 ;
        RECT 92.600 135.800 93.000 136.200 ;
        RECT 85.400 134.800 85.800 135.200 ;
        RECT 79.000 125.800 79.400 126.200 ;
        RECT 42.200 105.800 42.600 106.200 ;
        RECT 47.800 104.800 48.200 105.200 ;
        RECT 51.000 103.800 51.400 104.200 ;
        RECT 42.200 94.800 42.600 95.200 ;
        RECT 47.800 95.800 48.200 96.200 ;
        RECT 46.200 93.800 46.600 94.200 ;
        RECT 47.800 88.800 48.200 89.200 ;
        RECT 43.800 86.800 44.200 87.200 ;
        RECT 16.600 45.800 17.000 46.200 ;
        RECT 4.600 34.800 5.000 35.200 ;
        RECT 4.600 25.800 5.000 26.200 ;
        RECT 5.400 6.800 5.800 7.200 ;
        RECT 11.000 14.800 11.400 15.200 ;
        RECT 12.600 12.800 13.000 13.200 ;
        RECT 20.600 25.800 21.000 26.200 ;
        RECT 43.800 62.800 44.200 63.200 ;
        RECT 63.800 105.800 64.200 106.200 ;
        RECT 58.200 92.800 58.600 93.200 ;
        RECT 64.600 103.800 65.000 104.200 ;
        RECT 63.000 94.800 63.400 95.200 ;
        RECT 59.000 88.800 59.400 89.200 ;
        RECT 50.200 74.800 50.600 75.200 ;
        RECT 89.400 131.800 89.800 132.200 ;
        RECT 95.800 133.800 96.200 134.200 ;
        RECT 123.800 152.800 124.200 153.200 ;
        RECT 107.000 134.800 107.400 135.200 ;
        RECT 95.800 126.800 96.200 127.200 ;
        RECT 102.200 126.800 102.600 127.200 ;
        RECT 106.200 125.800 106.600 126.200 ;
        RECT 93.400 112.800 93.800 113.200 ;
        RECT 68.600 86.800 69.000 87.200 ;
        RECT 62.200 85.800 62.600 86.200 ;
        RECT 51.000 66.800 51.400 67.200 ;
        RECT 49.400 65.800 49.800 66.200 ;
        RECT 50.200 55.800 50.600 56.200 ;
        RECT 28.600 36.800 29.000 37.200 ;
        RECT 48.600 36.800 49.000 37.200 ;
        RECT 45.400 26.800 45.800 27.200 ;
        RECT 41.400 14.800 41.800 15.200 ;
        RECT 46.200 24.800 46.600 25.200 ;
        RECT 55.000 25.800 55.400 26.200 ;
        RECT 50.200 21.800 50.600 22.200 ;
        RECT 64.600 84.800 65.000 85.200 ;
        RECT 77.400 85.800 77.800 86.200 ;
        RECT 67.000 58.800 67.400 59.200 ;
        RECT 65.400 46.800 65.800 47.200 ;
        RECT 74.200 65.800 74.600 66.200 ;
        RECT 79.800 68.800 80.200 69.200 ;
        RECT 73.400 52.800 73.800 53.200 ;
        RECT 59.800 32.800 60.200 33.200 ;
        RECT 60.600 23.800 61.000 24.200 ;
        RECT 59.800 12.800 60.200 13.200 ;
        RECT 55.800 5.800 56.200 6.200 ;
        RECT 100.600 124.800 101.000 125.200 ;
        RECT 127.000 134.800 127.400 135.200 ;
        RECT 128.600 133.800 129.000 134.200 ;
        RECT 127.800 126.800 128.200 127.200 ;
        RECT 131.000 127.800 131.400 128.200 ;
        RECT 135.800 126.800 136.200 127.200 ;
        RECT 159.800 165.800 160.200 166.200 ;
        RECT 167.000 165.800 167.400 166.200 ;
        RECT 155.000 145.800 155.400 146.200 ;
        RECT 151.000 128.800 151.400 129.200 ;
        RECT 150.200 127.800 150.600 128.200 ;
        RECT 96.600 73.800 97.000 74.200 ;
        RECT 68.600 15.800 69.000 16.200 ;
        RECT 91.000 48.800 91.400 49.200 ;
        RECT 139.800 116.800 140.200 117.200 ;
        RECT 123.000 85.800 123.400 86.200 ;
        RECT 114.200 77.800 114.600 78.200 ;
        RECT 113.400 76.800 113.800 77.200 ;
        RECT 107.000 74.800 107.400 75.200 ;
        RECT 96.600 53.800 97.000 54.200 ;
        RECT 103.800 66.800 104.200 67.200 ;
        RECT 97.400 52.800 97.800 53.200 ;
        RECT 98.200 47.800 98.600 48.200 ;
        RECT 83.000 28.800 83.400 29.200 ;
        RECT 80.600 18.800 81.000 19.200 ;
        RECT 66.200 8.800 66.600 9.200 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 123.800 76.800 124.200 77.200 ;
        RECT 148.600 105.800 149.000 106.200 ;
        RECT 165.400 125.800 165.800 126.200 ;
        RECT 161.400 117.800 161.800 118.200 ;
        RECT 163.800 112.800 164.200 113.200 ;
        RECT 163.000 106.800 163.400 107.200 ;
        RECT 151.000 89.800 151.400 90.200 ;
        RECT 127.000 74.800 127.400 75.200 ;
        RECT 109.400 48.800 109.800 49.200 ;
        RECT 103.000 45.800 103.400 46.200 ;
        RECT 98.200 18.800 98.600 19.200 ;
        RECT 127.800 51.800 128.200 52.200 ;
        RECT 127.800 46.800 128.200 47.200 ;
        RECT 161.400 88.800 161.800 89.200 ;
        RECT 158.200 87.800 158.600 88.200 ;
        RECT 135.000 65.800 135.400 66.200 ;
        RECT 120.600 33.800 121.000 34.200 ;
        RECT 116.600 24.800 117.000 25.200 ;
        RECT 124.600 27.800 125.000 28.200 ;
        RECT 139.000 55.800 139.400 56.200 ;
        RECT 141.400 54.800 141.800 55.200 ;
        RECT 155.800 54.800 156.200 55.200 ;
        RECT 114.200 15.800 114.600 16.200 ;
        RECT 120.600 14.800 121.000 15.200 ;
        RECT 93.400 5.800 93.800 6.200 ;
        RECT 123.800 11.800 124.200 12.200 ;
        RECT 130.200 14.800 130.600 15.200 ;
        RECT 122.200 5.800 122.600 6.200 ;
        RECT 150.200 25.800 150.600 26.200 ;
        RECT 170.200 85.800 170.600 86.200 ;
        RECT 171.000 78.800 171.400 79.200 ;
        RECT 161.400 53.800 161.800 54.200 ;
        RECT 170.200 61.800 170.600 62.200 ;
        RECT 171.000 58.800 171.400 59.200 ;
        RECT 140.600 7.800 141.000 8.200 ;
        RECT 150.200 5.800 150.600 6.200 ;
        RECT 160.600 8.800 161.000 9.200 ;
        RECT 171.800 41.800 172.200 42.200 ;
        RECT 174.200 25.800 174.600 26.200 ;
        RECT 172.600 15.800 173.000 16.200 ;
        RECT 164.600 14.800 165.000 15.200 ;
      LAYER metal3 ;
        RECT 1.400 169.100 1.800 169.200 ;
        RECT 15.000 169.100 15.400 169.200 ;
        RECT 31.800 169.100 32.200 169.200 ;
        RECT 1.400 168.800 32.200 169.100 ;
        RECT 43.000 169.100 43.400 169.200 ;
        RECT 51.800 169.100 52.200 169.200 ;
        RECT 43.000 168.800 52.200 169.100 ;
        RECT 125.400 168.800 125.800 169.200 ;
        RECT 143.800 168.800 144.200 169.200 ;
        RECT 34.200 167.800 34.600 168.200 ;
        RECT 125.400 168.100 125.700 168.800 ;
        RECT 143.800 168.100 144.100 168.800 ;
        RECT 156.600 168.100 157.000 168.200 ;
        RECT 125.400 167.800 157.000 168.100 ;
        RECT 6.200 166.800 6.600 167.200 ;
        RECT 34.200 167.100 34.500 167.800 ;
        RECT 42.200 167.100 42.600 167.200 ;
        RECT 49.400 167.100 49.800 167.200 ;
        RECT 150.200 167.100 150.600 167.200 ;
        RECT 34.200 166.800 49.800 167.100 ;
        RECT 142.200 166.800 150.600 167.100 ;
        RECT 6.200 166.200 6.500 166.800 ;
        RECT 3.800 165.800 4.200 166.200 ;
        RECT 6.200 166.100 6.600 166.200 ;
        RECT 36.600 166.100 37.000 166.200 ;
        RECT 40.600 166.100 41.000 166.200 ;
        RECT 6.200 165.800 41.000 166.100 ;
        RECT 41.400 166.100 41.800 166.200 ;
        RECT 49.400 166.100 49.700 166.800 ;
        RECT 142.200 166.200 142.500 166.800 ;
        RECT 54.200 166.100 54.600 166.200 ;
        RECT 61.400 166.100 61.800 166.200 ;
        RECT 41.400 165.800 46.500 166.100 ;
        RECT 49.400 165.800 61.800 166.100 ;
        RECT 87.800 166.100 88.200 166.200 ;
        RECT 102.200 166.100 102.600 166.200 ;
        RECT 103.800 166.100 104.200 166.200 ;
        RECT 87.800 165.800 104.200 166.100 ;
        RECT 104.600 166.100 105.000 166.200 ;
        RECT 111.000 166.100 111.400 166.200 ;
        RECT 104.600 165.800 111.400 166.100 ;
        RECT 142.200 165.800 142.600 166.200 ;
        RECT 159.000 166.100 159.400 166.200 ;
        RECT 159.800 166.100 160.200 166.200 ;
        RECT 159.000 165.800 160.200 166.100 ;
        RECT 164.600 166.100 165.000 166.200 ;
        RECT 167.000 166.100 167.400 166.200 ;
        RECT 172.600 166.100 173.000 166.200 ;
        RECT 164.600 165.800 173.000 166.100 ;
        RECT 175.800 166.100 176.200 166.200 ;
        RECT 176.600 166.100 177.000 166.200 ;
        RECT 175.800 165.800 177.000 166.100 ;
        RECT 3.800 165.100 4.100 165.800 ;
        RECT 46.200 165.200 46.500 165.800 ;
        RECT 9.400 165.100 9.800 165.200 ;
        RECT 3.800 164.800 9.800 165.100 ;
        RECT 46.200 164.800 46.600 165.200 ;
        RECT 80.600 165.100 81.000 165.200 ;
        RECT 91.800 165.100 92.200 165.200 ;
        RECT 93.400 165.100 93.800 165.200 ;
        RECT 80.600 164.800 93.800 165.100 ;
        RECT 94.200 165.100 94.600 165.200 ;
        RECT 125.400 165.100 125.800 165.200 ;
        RECT 94.200 164.800 125.800 165.100 ;
        RECT 135.800 165.100 136.200 165.200 ;
        RECT 170.200 165.100 170.600 165.200 ;
        RECT 135.800 164.800 170.600 165.100 ;
        RECT 38.200 164.100 38.600 164.200 ;
        RECT 44.600 164.100 45.000 164.200 ;
        RECT 87.800 164.100 88.200 164.200 ;
        RECT 38.200 163.800 88.200 164.100 ;
        RECT 100.600 164.100 101.000 164.200 ;
        RECT 101.400 164.100 101.800 164.200 ;
        RECT 100.600 163.800 101.800 164.100 ;
        RECT 168.600 164.100 169.000 164.200 ;
        RECT 174.200 164.100 174.600 164.200 ;
        RECT 168.600 163.800 174.600 164.100 ;
        RECT 15.000 162.100 15.400 162.200 ;
        RECT 72.600 162.100 73.000 162.200 ;
        RECT 169.400 162.100 169.800 162.200 ;
        RECT 15.000 161.800 73.000 162.100 ;
        RECT 164.600 161.800 169.800 162.100 ;
        RECT 164.600 161.200 164.900 161.800 ;
        RECT 6.200 161.100 6.600 161.200 ;
        RECT 12.600 161.100 13.000 161.200 ;
        RECT 22.200 161.100 22.600 161.200 ;
        RECT 28.600 161.100 29.000 161.200 ;
        RECT 6.200 160.800 29.000 161.100 ;
        RECT 69.400 160.800 69.800 161.200 ;
        RECT 164.600 160.800 165.000 161.200 ;
        RECT 165.400 160.800 165.800 161.200 ;
        RECT 69.400 160.200 69.700 160.800 ;
        RECT 165.400 160.200 165.700 160.800 ;
        RECT 69.400 159.800 69.800 160.200 ;
        RECT 165.400 159.800 165.800 160.200 ;
        RECT 26.200 159.100 26.600 159.200 ;
        RECT 57.400 159.100 57.800 159.200 ;
        RECT 26.200 158.800 57.800 159.100 ;
        RECT 63.800 159.100 64.200 159.200 ;
        RECT 93.400 159.100 93.800 159.200 ;
        RECT 63.800 158.800 93.800 159.100 ;
        RECT 117.400 159.100 117.800 159.200 ;
        RECT 155.800 159.100 156.200 159.200 ;
        RECT 117.400 158.800 156.200 159.100 ;
        RECT 32.600 158.100 33.000 158.200 ;
        RECT 54.200 158.100 54.600 158.200 ;
        RECT 32.600 157.800 54.600 158.100 ;
        RECT 72.600 158.100 73.000 158.200 ;
        RECT 87.800 158.100 88.200 158.200 ;
        RECT 127.800 158.100 128.200 158.200 ;
        RECT 130.200 158.100 130.600 158.200 ;
        RECT 72.600 157.800 130.600 158.100 ;
        RECT 105.400 157.100 105.800 157.200 ;
        RECT 107.000 157.100 107.400 157.200 ;
        RECT 105.400 156.800 107.400 157.100 ;
        RECT 112.600 157.100 113.000 157.200 ;
        RECT 114.200 157.100 114.600 157.200 ;
        RECT 112.600 156.800 115.300 157.100 ;
        RECT 19.000 156.100 19.400 156.200 ;
        RECT 26.200 156.100 26.600 156.200 ;
        RECT 59.800 156.100 60.200 156.200 ;
        RECT 60.600 156.100 61.000 156.200 ;
        RECT 19.000 155.800 61.000 156.100 ;
        RECT 70.200 156.100 70.600 156.200 ;
        RECT 80.600 156.100 81.000 156.200 ;
        RECT 70.200 155.800 81.000 156.100 ;
        RECT 101.400 156.100 101.800 156.200 ;
        RECT 109.400 156.100 109.800 156.200 ;
        RECT 101.400 155.800 109.800 156.100 ;
        RECT 139.800 155.800 140.200 156.200 ;
        RECT 167.800 156.100 168.200 156.200 ;
        RECT 171.000 156.100 171.400 156.200 ;
        RECT 167.800 155.800 171.400 156.100 ;
        RECT 172.600 156.100 173.000 156.200 ;
        RECT 173.400 156.100 173.800 156.200 ;
        RECT 172.600 155.800 173.800 156.100 ;
        RECT 5.400 155.100 5.800 155.200 ;
        RECT 20.600 155.100 21.000 155.200 ;
        RECT 22.200 155.100 22.600 155.200 ;
        RECT 5.400 154.800 22.600 155.100 ;
        RECT 40.600 155.100 41.000 155.200 ;
        RECT 59.800 155.100 60.200 155.200 ;
        RECT 40.600 154.800 60.200 155.100 ;
        RECT 67.800 155.100 68.200 155.200 ;
        RECT 70.200 155.100 70.500 155.800 ;
        RECT 67.800 154.800 70.500 155.100 ;
        RECT 76.600 154.800 77.000 155.200 ;
        RECT 79.000 155.100 79.400 155.200 ;
        RECT 87.000 155.100 87.400 155.200 ;
        RECT 90.200 155.100 90.600 155.200 ;
        RECT 79.000 154.800 83.400 155.100 ;
        RECT 87.000 154.800 90.600 155.100 ;
        RECT 91.800 155.100 92.200 155.200 ;
        RECT 101.400 155.100 101.800 155.200 ;
        RECT 91.800 154.800 101.800 155.100 ;
        RECT 111.800 155.100 112.200 155.200 ;
        RECT 118.200 155.100 118.600 155.200 ;
        RECT 111.800 154.800 118.600 155.100 ;
        RECT 133.400 155.100 133.800 155.200 ;
        RECT 139.800 155.100 140.100 155.800 ;
        RECT 133.400 154.800 140.100 155.100 ;
        RECT 76.600 154.200 76.900 154.800 ;
        RECT 83.000 154.700 83.400 154.800 ;
        RECT 3.800 154.100 4.200 154.200 ;
        RECT 12.600 154.100 13.000 154.200 ;
        RECT 3.800 153.800 13.000 154.100 ;
        RECT 15.000 154.100 15.400 154.200 ;
        RECT 15.800 154.100 16.200 154.200 ;
        RECT 19.000 154.100 19.400 154.200 ;
        RECT 15.000 153.800 19.400 154.100 ;
        RECT 47.800 154.100 48.200 154.200 ;
        RECT 49.400 154.100 49.800 154.200 ;
        RECT 47.800 153.800 49.800 154.100 ;
        RECT 63.800 154.100 64.200 154.200 ;
        RECT 72.600 154.100 73.000 154.200 ;
        RECT 63.800 153.800 73.000 154.100 ;
        RECT 76.600 153.800 77.000 154.200 ;
        RECT 103.000 154.100 103.400 154.200 ;
        RECT 114.200 154.100 114.600 154.200 ;
        RECT 128.600 154.100 129.000 154.200 ;
        RECT 103.000 153.800 129.000 154.100 ;
        RECT 158.200 154.100 158.600 154.200 ;
        RECT 158.200 153.800 162.500 154.100 ;
        RECT 11.000 153.100 11.400 153.200 ;
        RECT 16.600 153.100 17.000 153.200 ;
        RECT 11.000 152.800 17.000 153.100 ;
        RECT 19.000 153.100 19.300 153.800 ;
        RECT 162.200 153.200 162.500 153.800 ;
        RECT 51.800 153.100 52.200 153.200 ;
        RECT 19.000 152.800 52.200 153.100 ;
        RECT 73.400 153.100 73.800 153.200 ;
        RECT 91.800 153.100 92.200 153.200 ;
        RECT 73.400 152.800 92.200 153.100 ;
        RECT 100.600 153.100 101.000 153.200 ;
        RECT 123.800 153.100 124.200 153.200 ;
        RECT 100.600 152.800 124.200 153.100 ;
        RECT 127.000 153.100 127.400 153.200 ;
        RECT 142.200 153.100 142.600 153.200 ;
        RECT 127.000 152.800 142.600 153.100 ;
        RECT 162.200 152.800 162.600 153.200 ;
        RECT 39.800 152.100 40.200 152.200 ;
        RECT 50.200 152.100 50.600 152.200 ;
        RECT 39.800 151.800 50.600 152.100 ;
        RECT 69.400 152.100 69.800 152.200 ;
        RECT 96.600 152.100 97.000 152.200 ;
        RECT 69.400 151.800 97.000 152.100 ;
        RECT 97.400 152.100 97.800 152.200 ;
        RECT 103.800 152.100 104.200 152.200 ;
        RECT 97.400 151.800 104.200 152.100 ;
        RECT 104.600 152.100 105.000 152.200 ;
        RECT 135.000 152.100 135.400 152.200 ;
        RECT 145.400 152.100 145.800 152.200 ;
        RECT 104.600 151.800 145.800 152.100 ;
        RECT 152.600 152.100 153.000 152.200 ;
        RECT 156.600 152.100 157.000 152.200 ;
        RECT 163.800 152.100 164.200 152.200 ;
        RECT 152.600 151.800 164.200 152.100 ;
        RECT 167.800 152.100 168.200 152.200 ;
        RECT 172.600 152.100 173.000 152.200 ;
        RECT 167.800 151.800 173.000 152.100 ;
        RECT 51.000 151.100 51.400 151.200 ;
        RECT 61.400 151.100 61.800 151.200 ;
        RECT 73.400 151.100 73.800 151.200 ;
        RECT 51.000 150.800 73.800 151.100 ;
        RECT 100.600 151.100 101.000 151.200 ;
        RECT 115.000 151.100 115.400 151.200 ;
        RECT 129.400 151.100 129.800 151.200 ;
        RECT 100.600 150.800 129.800 151.100 ;
        RECT 161.400 151.100 161.800 151.200 ;
        RECT 171.800 151.100 172.200 151.200 ;
        RECT 177.400 151.100 177.800 151.200 ;
        RECT 161.400 150.800 177.800 151.100 ;
        RECT 42.200 150.100 42.600 150.200 ;
        RECT 43.000 150.100 43.400 150.200 ;
        RECT 49.400 150.100 49.800 150.200 ;
        RECT 42.200 149.800 49.800 150.100 ;
        RECT 51.800 150.100 52.200 150.200 ;
        RECT 80.600 150.100 81.000 150.200 ;
        RECT 87.000 150.100 87.400 150.200 ;
        RECT 51.800 149.800 87.400 150.100 ;
        RECT 98.200 150.100 98.600 150.200 ;
        RECT 101.400 150.100 101.800 150.200 ;
        RECT 98.200 149.800 101.800 150.100 ;
        RECT 102.200 150.100 102.600 150.200 ;
        RECT 115.800 150.100 116.200 150.200 ;
        RECT 102.200 149.800 116.200 150.100 ;
        RECT 155.800 150.100 156.200 150.200 ;
        RECT 173.400 150.100 173.800 150.200 ;
        RECT 155.800 149.800 173.800 150.100 ;
        RECT 43.800 149.100 44.200 149.200 ;
        RECT 56.600 149.100 57.000 149.200 ;
        RECT 59.800 149.100 60.200 149.200 ;
        RECT 43.800 148.800 60.200 149.100 ;
        RECT 99.000 148.800 99.400 149.200 ;
        RECT 108.600 149.100 109.000 149.200 ;
        RECT 113.400 149.100 113.800 149.200 ;
        RECT 108.600 148.800 113.800 149.100 ;
        RECT 170.200 148.800 170.600 149.200 ;
        RECT 9.400 148.100 9.800 148.200 ;
        RECT 11.000 148.100 11.400 148.200 ;
        RECT 15.800 148.100 16.200 148.200 ;
        RECT 9.400 147.800 16.200 148.100 ;
        RECT 19.800 148.100 20.200 148.200 ;
        RECT 62.200 148.100 62.600 148.200 ;
        RECT 19.800 147.800 62.600 148.100 ;
        RECT 64.600 148.100 65.000 148.200 ;
        RECT 99.000 148.100 99.300 148.800 ;
        RECT 64.600 147.800 99.300 148.100 ;
        RECT 101.400 148.100 101.800 148.200 ;
        RECT 107.000 148.100 107.400 148.200 ;
        RECT 101.400 147.800 107.400 148.100 ;
        RECT 131.000 148.100 131.400 148.200 ;
        RECT 139.800 148.100 140.200 148.200 ;
        RECT 131.000 147.800 140.200 148.100 ;
        RECT 147.000 147.800 147.400 148.200 ;
        RECT 155.000 148.100 155.400 148.200 ;
        RECT 158.200 148.100 158.600 148.200 ;
        RECT 155.000 147.800 158.600 148.100 ;
        RECT 163.800 148.100 164.200 148.200 ;
        RECT 170.200 148.100 170.500 148.800 ;
        RECT 175.000 148.100 175.400 148.200 ;
        RECT 163.800 147.800 175.400 148.100 ;
        RECT 11.800 147.100 12.200 147.200 ;
        RECT 13.400 147.100 13.800 147.200 ;
        RECT 40.600 147.100 41.000 147.200 ;
        RECT 42.200 147.100 42.600 147.200 ;
        RECT 47.800 147.100 48.200 147.200 ;
        RECT 11.800 146.800 48.200 147.100 ;
        RECT 48.600 147.100 49.000 147.200 ;
        RECT 49.400 147.100 49.800 147.200 ;
        RECT 48.600 146.800 49.800 147.100 ;
        RECT 62.200 147.100 62.600 147.200 ;
        RECT 63.000 147.100 63.400 147.200 ;
        RECT 62.200 146.800 63.400 147.100 ;
        RECT 65.400 147.100 65.800 147.200 ;
        RECT 66.200 147.100 66.600 147.200 ;
        RECT 65.400 146.800 66.600 147.100 ;
        RECT 85.400 147.100 85.800 147.200 ;
        RECT 92.600 147.100 93.000 147.200 ;
        RECT 93.400 147.100 93.800 147.200 ;
        RECT 103.000 147.100 103.400 147.200 ;
        RECT 110.200 147.100 110.600 147.200 ;
        RECT 119.000 147.100 119.400 147.200 ;
        RECT 124.600 147.100 125.000 147.200 ;
        RECT 85.400 146.800 125.000 147.100 ;
        RECT 134.200 146.800 134.600 147.200 ;
        RECT 147.000 147.100 147.300 147.800 ;
        RECT 152.600 147.100 153.000 147.200 ;
        RECT 147.000 146.800 153.000 147.100 ;
        RECT 154.200 147.100 154.600 147.200 ;
        RECT 155.800 147.100 156.200 147.200 ;
        RECT 154.200 146.800 156.200 147.100 ;
        RECT 156.600 147.100 157.000 147.200 ;
        RECT 157.400 147.100 157.800 147.200 ;
        RECT 156.600 146.800 157.800 147.100 ;
        RECT 168.600 146.800 169.000 147.200 ;
        RECT 134.200 146.200 134.500 146.800 ;
        RECT 168.600 146.200 168.900 146.800 ;
        RECT 4.600 146.100 5.000 146.200 ;
        RECT 12.600 146.100 13.000 146.200 ;
        RECT 4.600 145.800 13.000 146.100 ;
        RECT 25.400 146.100 25.800 146.200 ;
        RECT 32.600 146.100 33.000 146.200 ;
        RECT 25.400 145.800 33.000 146.100 ;
        RECT 39.000 146.100 39.400 146.200 ;
        RECT 52.600 146.100 53.000 146.200 ;
        RECT 39.000 145.800 53.000 146.100 ;
        RECT 54.200 146.100 54.600 146.200 ;
        RECT 77.400 146.100 77.800 146.200 ;
        RECT 82.200 146.100 82.600 146.200 ;
        RECT 83.800 146.100 84.200 146.200 ;
        RECT 54.200 145.800 84.200 146.100 ;
        RECT 84.600 146.100 85.000 146.200 ;
        RECT 93.400 146.100 93.800 146.200 ;
        RECT 84.600 145.800 93.800 146.100 ;
        RECT 99.800 146.100 100.200 146.200 ;
        RECT 100.600 146.100 101.000 146.200 ;
        RECT 99.800 145.800 101.000 146.100 ;
        RECT 103.800 146.100 104.200 146.200 ;
        RECT 112.600 146.100 113.000 146.200 ;
        RECT 131.000 146.100 131.400 146.200 ;
        RECT 103.800 145.800 131.400 146.100 ;
        RECT 132.600 145.800 133.000 146.200 ;
        RECT 134.200 146.100 134.600 146.200 ;
        RECT 135.800 146.100 136.200 146.200 ;
        RECT 134.200 145.800 136.200 146.100 ;
        RECT 147.800 146.100 148.200 146.200 ;
        RECT 155.000 146.100 155.400 146.200 ;
        RECT 159.800 146.100 160.200 146.200 ;
        RECT 147.800 145.800 148.900 146.100 ;
        RECT 155.000 145.800 160.200 146.100 ;
        RECT 168.600 145.800 169.000 146.200 ;
        RECT 19.000 145.100 19.400 145.200 ;
        RECT 28.600 145.100 29.000 145.200 ;
        RECT 42.200 145.100 42.600 145.200 ;
        RECT 45.400 145.100 45.800 145.200 ;
        RECT 19.000 144.800 29.000 145.100 ;
        RECT 41.400 144.800 45.800 145.100 ;
        RECT 46.200 145.100 46.600 145.200 ;
        RECT 60.600 145.100 61.000 145.200 ;
        RECT 65.400 145.100 65.800 145.200 ;
        RECT 46.200 144.800 65.800 145.100 ;
        RECT 79.800 145.100 80.200 145.200 ;
        RECT 81.400 145.100 81.800 145.200 ;
        RECT 87.800 145.100 88.200 145.200 ;
        RECT 127.000 145.100 127.400 145.200 ;
        RECT 79.800 144.800 88.200 145.100 ;
        RECT 117.400 144.800 127.400 145.100 ;
        RECT 132.600 145.100 132.900 145.800 ;
        RECT 148.600 145.200 148.900 145.800 ;
        RECT 144.600 145.100 145.000 145.200 ;
        RECT 132.600 144.800 145.000 145.100 ;
        RECT 148.600 144.800 149.000 145.200 ;
        RECT 156.600 145.100 157.000 145.200 ;
        RECT 163.000 145.100 163.400 145.200 ;
        RECT 156.600 144.800 163.400 145.100 ;
        RECT 46.200 144.200 46.500 144.800 ;
        RECT 117.400 144.200 117.700 144.800 ;
        RECT 17.400 144.100 17.800 144.200 ;
        RECT 46.200 144.100 46.600 144.200 ;
        RECT 17.400 143.800 46.600 144.100 ;
        RECT 117.400 143.800 117.800 144.200 ;
        RECT 39.000 143.100 39.400 143.200 ;
        RECT 42.200 143.100 42.600 143.200 ;
        RECT 39.000 142.800 42.600 143.100 ;
        RECT 68.600 142.800 69.000 143.200 ;
        RECT 80.600 143.100 81.000 143.200 ;
        RECT 149.400 143.100 149.800 143.200 ;
        RECT 80.600 142.800 149.800 143.100 ;
        RECT 68.600 142.200 68.900 142.800 ;
        RECT 51.800 142.100 52.200 142.200 ;
        RECT 60.600 142.100 61.000 142.200 ;
        RECT 51.800 141.800 61.000 142.100 ;
        RECT 68.600 141.800 69.000 142.200 ;
        RECT 79.000 142.100 79.400 142.200 ;
        RECT 87.800 142.100 88.200 142.200 ;
        RECT 79.000 141.800 88.200 142.100 ;
        RECT 93.400 142.100 93.800 142.200 ;
        RECT 120.600 142.100 121.000 142.200 ;
        RECT 93.400 141.800 121.000 142.100 ;
        RECT 170.200 142.100 170.600 142.200 ;
        RECT 174.200 142.100 174.600 142.200 ;
        RECT 177.400 142.100 177.800 142.200 ;
        RECT 170.200 141.800 177.800 142.100 ;
        RECT 68.600 141.100 69.000 141.200 ;
        RECT 69.400 141.100 69.800 141.200 ;
        RECT 68.600 140.800 69.800 141.100 ;
        RECT 159.000 141.100 159.400 141.200 ;
        RECT 174.200 141.100 174.600 141.200 ;
        RECT 159.000 140.800 174.600 141.100 ;
        RECT 40.600 139.100 41.000 139.200 ;
        RECT 59.800 139.100 60.200 139.200 ;
        RECT 70.200 139.100 70.600 139.200 ;
        RECT 77.400 139.100 77.800 139.200 ;
        RECT 40.600 138.800 77.800 139.100 ;
        RECT 95.800 139.100 96.200 139.200 ;
        RECT 103.800 139.100 104.200 139.200 ;
        RECT 95.800 138.800 104.200 139.100 ;
        RECT 127.800 139.100 128.200 139.200 ;
        RECT 173.400 139.100 173.800 139.200 ;
        RECT 127.800 138.800 173.800 139.100 ;
        RECT 27.000 138.100 27.400 138.200 ;
        RECT 36.600 138.100 37.000 138.200 ;
        RECT 27.000 137.800 37.000 138.100 ;
        RECT 65.400 138.100 65.800 138.200 ;
        RECT 79.800 138.100 80.200 138.200 ;
        RECT 65.400 137.800 80.200 138.100 ;
        RECT 99.800 138.100 100.200 138.200 ;
        RECT 107.000 138.100 107.400 138.200 ;
        RECT 99.800 137.800 107.400 138.100 ;
        RECT 115.000 137.800 115.400 138.200 ;
        RECT 148.600 138.100 149.000 138.200 ;
        RECT 159.800 138.100 160.200 138.200 ;
        RECT 163.800 138.100 164.200 138.200 ;
        RECT 148.600 137.800 164.200 138.100 ;
        RECT 115.000 137.200 115.300 137.800 ;
        RECT 19.800 137.100 20.200 137.200 ;
        RECT 25.400 137.100 25.800 137.200 ;
        RECT 19.800 136.800 25.800 137.100 ;
        RECT 26.200 137.100 26.600 137.200 ;
        RECT 34.200 137.100 34.600 137.200 ;
        RECT 55.800 137.100 56.200 137.200 ;
        RECT 61.400 137.100 61.800 137.200 ;
        RECT 64.600 137.100 65.000 137.200 ;
        RECT 26.200 136.800 65.000 137.100 ;
        RECT 66.200 136.800 66.600 137.200 ;
        RECT 103.000 137.100 103.400 137.200 ;
        RECT 103.800 137.100 104.200 137.200 ;
        RECT 103.000 136.800 104.200 137.100 ;
        RECT 115.000 136.800 115.400 137.200 ;
        RECT 132.600 137.100 133.000 137.200 ;
        RECT 156.600 137.100 157.000 137.200 ;
        RECT 168.600 137.100 169.000 137.200 ;
        RECT 132.600 136.800 169.000 137.100 ;
        RECT 175.000 137.100 175.400 137.200 ;
        RECT 175.800 137.100 176.200 137.200 ;
        RECT 175.000 136.800 176.200 137.100 ;
        RECT 15.000 136.100 15.400 136.200 ;
        RECT 20.600 136.100 21.000 136.200 ;
        RECT 15.000 135.800 21.000 136.100 ;
        RECT 22.200 136.100 22.600 136.200 ;
        RECT 23.000 136.100 23.400 136.200 ;
        RECT 22.200 135.800 23.400 136.100 ;
        RECT 27.800 136.100 28.200 136.200 ;
        RECT 29.400 136.100 29.800 136.200 ;
        RECT 27.800 135.800 29.800 136.100 ;
        RECT 30.200 136.100 30.600 136.200 ;
        RECT 31.000 136.100 31.400 136.200 ;
        RECT 30.200 135.800 31.400 136.100 ;
        RECT 57.400 136.100 57.800 136.200 ;
        RECT 58.200 136.100 58.600 136.200 ;
        RECT 57.400 135.800 58.600 136.100 ;
        RECT 59.000 136.100 59.400 136.200 ;
        RECT 59.800 136.100 60.200 136.200 ;
        RECT 66.200 136.100 66.500 136.800 ;
        RECT 59.000 135.800 66.500 136.100 ;
        RECT 71.800 136.100 72.200 136.200 ;
        RECT 75.800 136.100 76.200 136.200 ;
        RECT 71.800 135.800 76.200 136.100 ;
        RECT 92.600 136.100 93.000 136.200 ;
        RECT 107.800 136.100 108.200 136.200 ;
        RECT 92.600 135.800 108.200 136.100 ;
        RECT 134.200 135.800 134.600 136.200 ;
        RECT 159.800 136.100 160.200 136.200 ;
        RECT 163.000 136.100 163.400 136.200 ;
        RECT 159.800 135.800 163.400 136.100 ;
        RECT 166.200 136.100 166.600 136.200 ;
        RECT 175.800 136.100 176.200 136.200 ;
        RECT 166.200 135.800 176.200 136.100 ;
        RECT 11.000 134.800 11.400 135.200 ;
        RECT 14.200 135.100 14.600 135.200 ;
        RECT 23.000 135.100 23.400 135.200 ;
        RECT 14.200 134.800 23.400 135.100 ;
        RECT 23.800 135.100 24.200 135.200 ;
        RECT 27.800 135.100 28.200 135.200 ;
        RECT 33.400 135.100 33.800 135.200 ;
        RECT 34.200 135.100 34.600 135.200 ;
        RECT 23.800 134.800 34.600 135.100 ;
        RECT 47.800 135.100 48.200 135.200 ;
        RECT 50.200 135.100 50.600 135.200 ;
        RECT 53.400 135.100 53.800 135.200 ;
        RECT 78.200 135.100 78.600 135.200 ;
        RECT 47.800 134.800 78.600 135.100 ;
        RECT 85.400 135.100 85.800 135.200 ;
        RECT 87.000 135.100 87.400 135.200 ;
        RECT 85.400 134.800 87.400 135.100 ;
        RECT 92.600 135.100 93.000 135.200 ;
        RECT 104.600 135.100 105.000 135.200 ;
        RECT 107.000 135.100 107.400 135.200 ;
        RECT 92.600 134.800 107.400 135.100 ;
        RECT 113.400 135.100 113.800 135.200 ;
        RECT 114.200 135.100 114.600 135.200 ;
        RECT 127.000 135.100 127.400 135.200 ;
        RECT 130.200 135.100 130.600 135.200 ;
        RECT 113.400 134.800 116.100 135.100 ;
        RECT 127.000 134.800 130.600 135.100 ;
        RECT 134.200 135.100 134.500 135.800 ;
        RECT 143.800 135.100 144.200 135.200 ;
        RECT 134.200 134.800 144.200 135.100 ;
        RECT 157.400 134.800 157.800 135.200 ;
        RECT 159.000 135.100 159.400 135.200 ;
        RECT 165.400 135.100 165.800 135.200 ;
        RECT 167.000 135.100 167.400 135.200 ;
        RECT 159.000 134.800 167.400 135.100 ;
        RECT 171.000 135.100 171.400 135.200 ;
        RECT 178.200 135.100 178.600 135.200 ;
        RECT 171.000 134.800 178.600 135.100 ;
        RECT 6.200 134.100 6.600 134.200 ;
        RECT 11.000 134.100 11.300 134.800 ;
        RECT 115.800 134.200 116.100 134.800 ;
        RECT 157.400 134.200 157.700 134.800 ;
        RECT 6.200 133.800 11.300 134.100 ;
        RECT 31.000 134.100 31.400 134.200 ;
        RECT 35.800 134.100 36.200 134.200 ;
        RECT 31.000 133.800 36.200 134.100 ;
        RECT 51.800 134.100 52.200 134.200 ;
        RECT 53.400 134.100 53.800 134.200 ;
        RECT 51.800 133.800 53.800 134.100 ;
        RECT 55.800 134.100 56.200 134.200 ;
        RECT 56.600 134.100 57.000 134.200 ;
        RECT 55.800 133.800 57.000 134.100 ;
        RECT 63.800 134.100 64.200 134.200 ;
        RECT 72.600 134.100 73.000 134.200 ;
        RECT 63.800 133.800 73.000 134.100 ;
        RECT 95.000 134.100 95.400 134.200 ;
        RECT 95.800 134.100 96.200 134.200 ;
        RECT 95.000 133.800 96.200 134.100 ;
        RECT 102.200 134.100 102.600 134.200 ;
        RECT 103.000 134.100 103.400 134.200 ;
        RECT 102.200 133.800 103.400 134.100 ;
        RECT 115.800 133.800 116.200 134.200 ;
        RECT 119.800 134.100 120.200 134.200 ;
        RECT 128.600 134.100 129.000 134.200 ;
        RECT 119.800 133.800 129.000 134.100 ;
        RECT 147.000 134.100 147.400 134.200 ;
        RECT 153.400 134.100 153.800 134.200 ;
        RECT 147.000 133.800 153.800 134.100 ;
        RECT 157.400 134.100 157.800 134.200 ;
        RECT 172.600 134.100 173.000 134.200 ;
        RECT 157.400 133.800 173.000 134.100 ;
        RECT 39.000 133.100 39.400 133.200 ;
        RECT 41.400 133.100 41.800 133.200 ;
        RECT 39.000 132.800 41.800 133.100 ;
        RECT 43.000 133.100 43.400 133.200 ;
        RECT 52.600 133.100 53.000 133.200 ;
        RECT 43.000 132.800 53.000 133.100 ;
        RECT 56.600 133.100 56.900 133.800 ;
        RECT 61.400 133.100 61.800 133.200 ;
        RECT 56.600 132.800 61.800 133.100 ;
        RECT 67.800 133.100 68.200 133.200 ;
        RECT 71.000 133.100 71.400 133.200 ;
        RECT 67.800 132.800 71.400 133.100 ;
        RECT 82.200 133.100 82.600 133.200 ;
        RECT 83.000 133.100 83.400 133.200 ;
        RECT 82.200 132.800 83.400 133.100 ;
        RECT 95.800 133.100 96.100 133.800 ;
        RECT 101.400 133.100 101.800 133.200 ;
        RECT 108.600 133.100 109.000 133.200 ;
        RECT 95.800 132.800 109.000 133.100 ;
        RECT 119.000 133.100 119.400 133.200 ;
        RECT 123.800 133.100 124.200 133.200 ;
        RECT 119.000 132.800 124.200 133.100 ;
        RECT 131.800 133.100 132.200 133.200 ;
        RECT 132.600 133.100 133.000 133.200 ;
        RECT 135.000 133.100 135.400 133.200 ;
        RECT 131.800 132.800 135.400 133.100 ;
        RECT 143.000 133.100 143.400 133.200 ;
        RECT 154.200 133.100 154.600 133.200 ;
        RECT 143.000 132.800 154.600 133.100 ;
        RECT 159.800 132.800 160.200 133.200 ;
        RECT 166.200 133.100 166.600 133.200 ;
        RECT 167.000 133.100 167.400 133.200 ;
        RECT 166.200 132.800 167.400 133.100 ;
        RECT 167.800 133.100 168.200 133.200 ;
        RECT 168.600 133.100 169.000 133.200 ;
        RECT 167.800 132.800 169.000 133.100 ;
        RECT 169.400 133.100 169.800 133.200 ;
        RECT 178.200 133.100 178.600 133.200 ;
        RECT 169.400 132.800 178.600 133.100 ;
        RECT 159.800 132.200 160.100 132.800 ;
        RECT 4.600 132.100 5.000 132.200 ;
        RECT 6.200 132.100 6.600 132.200 ;
        RECT 19.800 132.100 20.200 132.200 ;
        RECT 37.400 132.100 37.800 132.200 ;
        RECT 4.600 131.800 37.800 132.100 ;
        RECT 44.600 131.800 45.000 132.200 ;
        RECT 49.400 132.100 49.800 132.200 ;
        RECT 58.200 132.100 58.600 132.200 ;
        RECT 49.400 131.800 58.600 132.100 ;
        RECT 73.400 131.800 73.800 132.200 ;
        RECT 83.000 132.100 83.400 132.200 ;
        RECT 87.800 132.100 88.200 132.200 ;
        RECT 83.000 131.800 88.200 132.100 ;
        RECT 89.400 132.100 89.800 132.200 ;
        RECT 140.600 132.100 141.000 132.200 ;
        RECT 89.400 131.800 141.000 132.100 ;
        RECT 147.800 131.800 148.200 132.200 ;
        RECT 159.800 131.800 160.200 132.200 ;
        RECT 167.000 132.100 167.400 132.200 ;
        RECT 171.000 132.100 171.400 132.200 ;
        RECT 167.000 131.800 171.400 132.100 ;
        RECT 44.600 131.200 44.900 131.800 ;
        RECT 73.400 131.200 73.700 131.800 ;
        RECT 147.800 131.200 148.100 131.800 ;
        RECT 6.200 131.100 6.600 131.200 ;
        RECT 9.400 131.100 9.800 131.200 ;
        RECT 23.000 131.100 23.400 131.200 ;
        RECT 6.200 130.800 23.400 131.100 ;
        RECT 44.600 130.800 45.000 131.200 ;
        RECT 45.400 130.800 45.800 131.200 ;
        RECT 73.400 130.800 73.800 131.200 ;
        RECT 81.400 131.100 81.800 131.200 ;
        RECT 83.800 131.100 84.200 131.200 ;
        RECT 81.400 130.800 84.200 131.100 ;
        RECT 103.800 130.800 104.200 131.200 ;
        RECT 115.000 131.100 115.400 131.200 ;
        RECT 129.400 131.100 129.800 131.200 ;
        RECT 115.000 130.800 129.800 131.100 ;
        RECT 147.800 130.800 148.200 131.200 ;
        RECT 151.000 131.100 151.400 131.200 ;
        RECT 166.200 131.100 166.600 131.200 ;
        RECT 151.000 130.800 166.600 131.100 ;
        RECT 45.400 130.200 45.700 130.800 ;
        RECT 103.800 130.200 104.100 130.800 ;
        RECT 45.400 129.800 45.800 130.200 ;
        RECT 51.000 130.100 51.400 130.200 ;
        RECT 59.000 130.100 59.400 130.200 ;
        RECT 63.800 130.100 64.200 130.200 ;
        RECT 51.000 129.800 64.200 130.100 ;
        RECT 67.000 130.100 67.400 130.200 ;
        RECT 70.200 130.100 70.600 130.200 ;
        RECT 67.000 129.800 70.600 130.100 ;
        RECT 103.800 129.800 104.200 130.200 ;
        RECT 107.800 130.100 108.200 130.200 ;
        RECT 110.200 130.100 110.600 130.200 ;
        RECT 107.800 129.800 110.600 130.100 ;
        RECT 131.000 130.100 131.400 130.200 ;
        RECT 160.600 130.100 161.000 130.200 ;
        RECT 131.000 129.800 161.000 130.100 ;
        RECT 35.800 129.100 36.200 129.200 ;
        RECT 43.000 129.100 43.400 129.200 ;
        RECT 63.000 129.100 63.400 129.200 ;
        RECT 75.800 129.100 76.200 129.200 ;
        RECT 35.800 128.800 63.400 129.100 ;
        RECT 67.800 128.800 76.200 129.100 ;
        RECT 107.000 129.100 107.400 129.200 ;
        RECT 116.600 129.100 117.000 129.200 ;
        RECT 127.000 129.100 127.400 129.200 ;
        RECT 107.000 128.800 127.400 129.100 ;
        RECT 151.000 129.100 151.400 129.200 ;
        RECT 151.800 129.100 152.200 129.200 ;
        RECT 151.000 128.800 152.200 129.100 ;
        RECT 11.800 128.100 12.200 128.200 ;
        RECT 22.200 128.100 22.600 128.200 ;
        RECT 11.800 127.800 22.600 128.100 ;
        RECT 35.000 128.100 35.400 128.200 ;
        RECT 53.400 128.100 53.800 128.200 ;
        RECT 67.800 128.100 68.100 128.800 ;
        RECT 35.000 127.800 53.800 128.100 ;
        RECT 60.600 127.800 68.100 128.100 ;
        RECT 68.600 127.800 69.000 128.200 ;
        RECT 85.400 127.800 85.800 128.200 ;
        RECT 96.600 128.100 97.000 128.200 ;
        RECT 106.200 128.100 106.600 128.200 ;
        RECT 96.600 127.800 106.600 128.100 ;
        RECT 115.800 127.800 116.200 128.200 ;
        RECT 131.000 128.100 131.400 128.200 ;
        RECT 123.800 127.800 131.400 128.100 ;
        RECT 134.200 127.800 134.600 128.200 ;
        RECT 149.400 128.100 149.800 128.200 ;
        RECT 150.200 128.100 150.600 128.200 ;
        RECT 149.400 127.800 150.600 128.100 ;
        RECT 163.000 128.100 163.400 128.200 ;
        RECT 164.600 128.100 165.000 128.200 ;
        RECT 163.000 127.800 165.000 128.100 ;
        RECT 167.000 128.100 167.400 128.200 ;
        RECT 173.400 128.100 173.800 128.200 ;
        RECT 167.000 127.800 173.800 128.100 ;
        RECT 176.600 127.800 177.000 128.200 ;
        RECT 60.600 127.200 60.900 127.800 ;
        RECT 68.600 127.200 68.900 127.800 ;
        RECT 85.400 127.200 85.700 127.800 ;
        RECT 29.400 127.100 29.800 127.200 ;
        RECT 39.000 127.100 39.400 127.200 ;
        RECT 29.400 126.800 39.400 127.100 ;
        RECT 43.800 127.100 44.200 127.200 ;
        RECT 45.400 127.100 45.800 127.200 ;
        RECT 43.800 126.800 45.800 127.100 ;
        RECT 52.600 127.100 53.000 127.200 ;
        RECT 53.400 127.100 53.800 127.200 ;
        RECT 52.600 126.800 53.800 127.100 ;
        RECT 60.600 126.800 61.000 127.200 ;
        RECT 61.400 127.100 61.800 127.200 ;
        RECT 63.800 127.100 64.200 127.200 ;
        RECT 67.800 127.100 68.200 127.200 ;
        RECT 61.400 126.800 68.200 127.100 ;
        RECT 68.600 126.800 69.000 127.200 ;
        RECT 85.400 126.800 85.800 127.200 ;
        RECT 86.200 127.100 86.600 127.200 ;
        RECT 95.800 127.100 96.200 127.200 ;
        RECT 86.200 126.800 96.200 127.100 ;
        RECT 101.400 127.100 101.800 127.200 ;
        RECT 102.200 127.100 102.600 127.200 ;
        RECT 101.400 126.800 102.600 127.100 ;
        RECT 115.800 127.100 116.100 127.800 ;
        RECT 123.800 127.200 124.100 127.800 ;
        RECT 134.200 127.200 134.500 127.800 ;
        RECT 176.600 127.200 176.900 127.800 ;
        RECT 120.600 127.100 121.000 127.200 ;
        RECT 115.800 126.800 121.000 127.100 ;
        RECT 123.800 126.800 124.200 127.200 ;
        RECT 127.800 127.100 128.200 127.200 ;
        RECT 131.800 127.100 132.200 127.200 ;
        RECT 127.800 126.800 132.200 127.100 ;
        RECT 134.200 126.800 134.600 127.200 ;
        RECT 135.800 127.100 136.200 127.200 ;
        RECT 147.000 127.100 147.400 127.200 ;
        RECT 135.000 126.800 147.400 127.100 ;
        RECT 163.800 127.100 164.200 127.200 ;
        RECT 168.600 127.100 169.000 127.200 ;
        RECT 163.800 126.800 169.000 127.100 ;
        RECT 176.600 126.800 177.000 127.200 ;
        RECT 2.200 126.100 2.600 126.200 ;
        RECT 5.400 126.100 5.800 126.200 ;
        RECT 2.200 125.800 5.800 126.100 ;
        RECT 11.000 126.100 11.400 126.200 ;
        RECT 39.000 126.100 39.400 126.200 ;
        RECT 54.200 126.100 54.600 126.200 ;
        RECT 11.000 125.800 16.100 126.100 ;
        RECT 39.000 125.800 54.600 126.100 ;
        RECT 59.800 126.100 60.200 126.200 ;
        RECT 60.600 126.100 61.000 126.200 ;
        RECT 66.200 126.100 66.600 126.200 ;
        RECT 72.600 126.100 73.000 126.200 ;
        RECT 59.800 125.800 61.000 126.100 ;
        RECT 65.400 125.800 73.000 126.100 ;
        RECT 79.000 126.100 79.400 126.200 ;
        RECT 99.800 126.100 100.200 126.200 ;
        RECT 79.000 125.800 100.200 126.100 ;
        RECT 103.000 126.100 103.400 126.200 ;
        RECT 106.200 126.100 106.600 126.200 ;
        RECT 137.400 126.100 137.800 126.200 ;
        RECT 103.000 125.800 137.800 126.100 ;
        RECT 165.400 125.800 165.800 126.200 ;
        RECT 166.200 125.800 166.600 126.200 ;
        RECT 168.600 126.100 168.900 126.800 ;
        RECT 171.800 126.100 172.200 126.200 ;
        RECT 168.600 125.800 172.200 126.100 ;
        RECT 15.800 125.200 16.100 125.800 ;
        RECT 165.400 125.200 165.700 125.800 ;
        RECT 3.800 125.100 4.200 125.200 ;
        RECT 10.200 125.100 10.600 125.200 ;
        RECT 3.800 124.800 10.600 125.100 ;
        RECT 15.800 124.800 16.200 125.200 ;
        RECT 21.400 125.100 21.800 125.200 ;
        RECT 28.600 125.100 29.000 125.200 ;
        RECT 43.800 125.100 44.200 125.200 ;
        RECT 63.800 125.100 64.200 125.200 ;
        RECT 21.400 124.800 64.200 125.100 ;
        RECT 64.600 125.100 65.000 125.200 ;
        RECT 71.800 125.100 72.200 125.200 ;
        RECT 64.600 124.800 72.200 125.100 ;
        RECT 74.200 125.100 74.600 125.200 ;
        RECT 77.400 125.100 77.800 125.200 ;
        RECT 74.200 124.800 77.800 125.100 ;
        RECT 99.800 125.100 100.200 125.200 ;
        RECT 100.600 125.100 101.000 125.200 ;
        RECT 99.800 124.800 101.000 125.100 ;
        RECT 103.800 125.100 104.200 125.200 ;
        RECT 135.800 125.100 136.200 125.200 ;
        RECT 161.400 125.100 161.800 125.200 ;
        RECT 162.200 125.100 162.600 125.200 ;
        RECT 103.800 124.800 162.600 125.100 ;
        RECT 165.400 124.800 165.800 125.200 ;
        RECT 166.200 125.100 166.500 125.800 ;
        RECT 173.400 125.100 173.800 125.200 ;
        RECT 166.200 124.800 173.800 125.100 ;
        RECT 4.600 124.100 5.000 124.200 ;
        RECT 15.800 124.100 16.200 124.200 ;
        RECT 4.600 123.800 16.200 124.100 ;
        RECT 25.400 124.100 25.800 124.200 ;
        RECT 39.800 124.100 40.200 124.200 ;
        RECT 25.400 123.800 40.200 124.100 ;
        RECT 63.800 124.100 64.200 124.200 ;
        RECT 64.600 124.100 65.000 124.200 ;
        RECT 66.200 124.100 66.600 124.200 ;
        RECT 63.800 123.800 66.600 124.100 ;
        RECT 72.600 124.100 73.000 124.200 ;
        RECT 102.200 124.100 102.600 124.200 ;
        RECT 114.200 124.100 114.600 124.200 ;
        RECT 72.600 123.800 114.600 124.100 ;
        RECT 133.400 124.100 133.800 124.200 ;
        RECT 159.800 124.100 160.200 124.200 ;
        RECT 133.400 123.800 160.200 124.100 ;
        RECT 170.200 124.100 170.600 124.200 ;
        RECT 179.800 124.100 180.200 124.200 ;
        RECT 170.200 123.800 180.200 124.100 ;
        RECT 39.800 123.100 40.200 123.200 ;
        RECT 60.600 123.100 61.000 123.200 ;
        RECT 39.800 122.800 61.000 123.100 ;
        RECT 72.600 123.100 73.000 123.200 ;
        RECT 99.000 123.100 99.400 123.200 ;
        RECT 115.000 123.100 115.400 123.200 ;
        RECT 128.600 123.100 129.000 123.200 ;
        RECT 72.600 122.800 129.000 123.100 ;
        RECT 129.400 123.100 129.800 123.200 ;
        RECT 133.400 123.100 133.800 123.200 ;
        RECT 129.400 122.800 133.800 123.100 ;
        RECT 37.400 122.100 37.800 122.200 ;
        RECT 41.400 122.100 41.800 122.200 ;
        RECT 37.400 121.800 41.800 122.100 ;
        RECT 51.800 122.100 52.200 122.200 ;
        RECT 76.600 122.100 77.000 122.200 ;
        RECT 51.800 121.800 77.000 122.100 ;
        RECT 140.600 122.100 141.000 122.200 ;
        RECT 175.000 122.100 175.400 122.200 ;
        RECT 140.600 121.800 175.400 122.100 ;
        RECT 179.800 121.800 180.200 122.200 ;
        RECT 179.800 121.200 180.100 121.800 ;
        RECT 96.600 121.100 97.000 121.200 ;
        RECT 97.400 121.100 97.800 121.200 ;
        RECT 96.600 120.800 97.800 121.100 ;
        RECT 162.200 121.100 162.600 121.200 ;
        RECT 167.000 121.100 167.400 121.200 ;
        RECT 162.200 120.800 167.400 121.100 ;
        RECT 179.800 120.800 180.200 121.200 ;
        RECT 7.000 119.100 7.400 119.200 ;
        RECT 7.000 118.800 28.900 119.100 ;
        RECT 25.400 117.800 25.800 118.200 ;
        RECT 28.600 118.100 28.900 118.800 ;
        RECT 95.800 118.800 96.200 119.200 ;
        RECT 39.800 118.100 40.200 118.200 ;
        RECT 28.600 117.800 40.200 118.100 ;
        RECT 95.800 118.100 96.100 118.800 ;
        RECT 97.400 118.100 97.800 118.200 ;
        RECT 95.800 117.800 97.800 118.100 ;
        RECT 161.400 118.100 161.800 118.200 ;
        RECT 167.000 118.100 167.400 118.200 ;
        RECT 161.400 117.800 167.400 118.100 ;
        RECT 169.400 118.100 169.800 118.200 ;
        RECT 171.800 118.100 172.200 118.200 ;
        RECT 169.400 117.800 172.200 118.100 ;
        RECT 25.400 117.200 25.700 117.800 ;
        RECT 2.200 117.100 2.600 117.200 ;
        RECT 9.400 117.100 9.800 117.200 ;
        RECT 2.200 116.800 9.800 117.100 ;
        RECT 25.400 116.800 25.800 117.200 ;
        RECT 43.000 117.100 43.400 117.200 ;
        RECT 50.200 117.100 50.600 117.200 ;
        RECT 43.000 116.800 50.600 117.100 ;
        RECT 71.800 117.100 72.200 117.200 ;
        RECT 74.200 117.100 74.600 117.200 ;
        RECT 71.800 116.800 74.600 117.100 ;
        RECT 83.000 117.100 83.400 117.200 ;
        RECT 94.200 117.100 94.600 117.200 ;
        RECT 83.000 116.800 94.600 117.100 ;
        RECT 95.000 117.100 95.400 117.200 ;
        RECT 95.800 117.100 96.200 117.200 ;
        RECT 95.000 116.800 96.200 117.100 ;
        RECT 96.600 117.100 97.000 117.200 ;
        RECT 99.000 117.100 99.400 117.200 ;
        RECT 96.600 116.800 99.400 117.100 ;
        RECT 112.600 116.800 113.000 117.200 ;
        RECT 139.800 117.100 140.200 117.200 ;
        RECT 171.000 117.100 171.400 117.200 ;
        RECT 139.800 116.800 171.400 117.100 ;
        RECT 3.800 116.100 4.200 116.200 ;
        RECT 7.800 116.100 8.200 116.200 ;
        RECT 16.600 116.100 17.000 116.200 ;
        RECT 31.800 116.100 32.200 116.200 ;
        RECT 44.600 116.100 45.000 116.200 ;
        RECT 47.800 116.100 48.200 116.200 ;
        RECT 3.800 115.800 48.200 116.100 ;
        RECT 63.800 116.100 64.200 116.200 ;
        RECT 92.600 116.100 93.000 116.200 ;
        RECT 63.800 115.800 93.000 116.100 ;
        RECT 112.600 116.100 112.900 116.800 ;
        RECT 121.400 116.100 121.800 116.200 ;
        RECT 112.600 115.800 121.800 116.100 ;
        RECT 132.600 116.100 133.000 116.200 ;
        RECT 157.400 116.100 157.800 116.200 ;
        RECT 132.600 115.800 157.800 116.100 ;
        RECT 159.800 116.100 160.200 116.200 ;
        RECT 165.400 116.100 165.800 116.200 ;
        RECT 159.800 115.800 165.800 116.100 ;
        RECT 169.400 115.800 169.800 116.200 ;
        RECT 169.400 115.200 169.700 115.800 ;
        RECT 2.200 115.100 2.600 115.200 ;
        RECT 5.400 115.100 5.800 115.200 ;
        RECT 2.200 114.800 5.800 115.100 ;
        RECT 15.800 115.100 16.200 115.200 ;
        RECT 36.600 115.100 37.000 115.200 ;
        RECT 15.800 114.800 37.000 115.100 ;
        RECT 47.000 115.100 47.400 115.200 ;
        RECT 56.600 115.100 57.000 115.200 ;
        RECT 47.000 114.800 57.000 115.100 ;
        RECT 71.000 115.100 71.400 115.200 ;
        RECT 72.600 115.100 73.000 115.200 ;
        RECT 71.000 114.800 73.000 115.100 ;
        RECT 75.000 115.100 75.400 115.200 ;
        RECT 78.200 115.100 78.600 115.200 ;
        RECT 75.000 114.800 78.600 115.100 ;
        RECT 84.600 115.100 85.000 115.200 ;
        RECT 85.400 115.100 85.800 115.200 ;
        RECT 84.600 114.800 85.800 115.100 ;
        RECT 91.000 115.100 91.400 115.200 ;
        RECT 104.600 115.100 105.000 115.200 ;
        RECT 91.000 114.800 105.000 115.100 ;
        RECT 115.000 115.100 115.400 115.200 ;
        RECT 160.600 115.100 161.000 115.200 ;
        RECT 115.000 114.800 161.000 115.100 ;
        RECT 169.400 114.800 169.800 115.200 ;
        RECT 115.000 114.200 115.300 114.800 ;
        RECT 6.200 113.800 6.600 114.200 ;
        RECT 18.200 114.100 18.600 114.200 ;
        RECT 19.800 114.100 20.200 114.200 ;
        RECT 18.200 113.800 20.200 114.100 ;
        RECT 32.600 114.100 33.000 114.200 ;
        RECT 35.000 114.100 35.400 114.200 ;
        RECT 32.600 113.800 35.400 114.100 ;
        RECT 42.200 114.100 42.600 114.200 ;
        RECT 86.200 114.100 86.600 114.200 ;
        RECT 98.200 114.100 98.600 114.200 ;
        RECT 107.000 114.100 107.400 114.200 ;
        RECT 42.200 113.800 107.400 114.100 ;
        RECT 115.000 113.800 115.400 114.200 ;
        RECT 135.800 114.100 136.200 114.200 ;
        RECT 146.200 114.100 146.600 114.200 ;
        RECT 135.800 113.800 146.600 114.100 ;
        RECT 159.800 114.100 160.200 114.200 ;
        RECT 161.400 114.100 161.800 114.200 ;
        RECT 159.800 113.800 161.800 114.100 ;
        RECT 162.200 114.100 162.600 114.200 ;
        RECT 163.000 114.100 163.400 114.200 ;
        RECT 162.200 113.800 163.400 114.100 ;
        RECT 166.200 114.100 166.600 114.200 ;
        RECT 170.200 114.100 170.600 114.200 ;
        RECT 166.200 113.800 170.600 114.100 ;
        RECT 6.200 113.100 6.500 113.800 ;
        RECT 15.800 113.100 16.200 113.200 ;
        RECT 6.200 112.800 16.200 113.100 ;
        RECT 25.400 113.100 25.800 113.200 ;
        RECT 34.200 113.100 34.600 113.200 ;
        RECT 25.400 112.800 34.600 113.100 ;
        RECT 35.000 113.100 35.400 113.200 ;
        RECT 42.200 113.100 42.600 113.200 ;
        RECT 35.000 112.800 42.600 113.100 ;
        RECT 65.400 113.100 65.800 113.200 ;
        RECT 69.400 113.100 69.800 113.200 ;
        RECT 65.400 112.800 69.800 113.100 ;
        RECT 75.800 113.100 76.200 113.200 ;
        RECT 83.000 113.100 83.400 113.200 ;
        RECT 75.800 112.800 83.400 113.100 ;
        RECT 93.400 113.100 93.800 113.200 ;
        RECT 96.600 113.100 97.000 113.200 ;
        RECT 93.400 112.800 97.000 113.100 ;
        RECT 107.800 113.100 108.200 113.200 ;
        RECT 121.400 113.100 121.800 113.200 ;
        RECT 107.800 112.800 121.800 113.100 ;
        RECT 135.800 113.100 136.200 113.200 ;
        RECT 143.800 113.100 144.200 113.200 ;
        RECT 144.600 113.100 145.000 113.200 ;
        RECT 152.600 113.100 153.000 113.200 ;
        RECT 135.800 112.800 153.000 113.100 ;
        RECT 155.000 113.100 155.400 113.200 ;
        RECT 163.800 113.100 164.200 113.200 ;
        RECT 155.000 112.800 164.200 113.100 ;
        RECT 164.600 113.100 165.000 113.200 ;
        RECT 173.400 113.100 173.800 113.200 ;
        RECT 164.600 112.800 173.800 113.100 ;
        RECT 23.000 112.100 23.400 112.200 ;
        RECT 31.000 112.100 31.400 112.200 ;
        RECT 23.000 111.800 31.400 112.100 ;
        RECT 36.600 112.100 37.000 112.200 ;
        RECT 47.000 112.100 47.400 112.200 ;
        RECT 36.600 111.800 47.400 112.100 ;
        RECT 81.400 112.100 81.800 112.200 ;
        RECT 87.800 112.100 88.200 112.200 ;
        RECT 81.400 111.800 88.200 112.100 ;
        RECT 101.400 112.100 101.800 112.200 ;
        RECT 109.400 112.100 109.800 112.200 ;
        RECT 115.000 112.100 115.400 112.200 ;
        RECT 101.400 111.800 115.400 112.100 ;
        RECT 137.400 112.100 137.800 112.200 ;
        RECT 147.000 112.100 147.400 112.200 ;
        RECT 137.400 111.800 147.400 112.100 ;
        RECT 151.000 112.100 151.400 112.200 ;
        RECT 151.800 112.100 152.200 112.200 ;
        RECT 151.000 111.800 152.200 112.100 ;
        RECT 31.000 111.100 31.400 111.200 ;
        RECT 36.600 111.100 36.900 111.800 ;
        RECT 31.000 110.800 36.900 111.100 ;
        RECT 59.800 111.100 60.200 111.200 ;
        RECT 63.000 111.100 63.400 111.200 ;
        RECT 59.800 110.800 63.400 111.100 ;
        RECT 99.000 111.100 99.400 111.200 ;
        RECT 107.000 111.100 107.400 111.200 ;
        RECT 99.000 110.800 107.400 111.100 ;
        RECT 172.600 111.100 173.000 111.200 ;
        RECT 174.200 111.100 174.600 111.200 ;
        RECT 172.600 110.800 174.600 111.100 ;
        RECT 54.200 110.100 54.600 110.200 ;
        RECT 80.600 110.100 81.000 110.200 ;
        RECT 54.200 109.800 81.000 110.100 ;
        RECT 96.600 110.100 97.000 110.200 ;
        RECT 99.000 110.100 99.400 110.200 ;
        RECT 96.600 109.800 99.400 110.100 ;
        RECT 157.400 110.100 157.800 110.200 ;
        RECT 162.200 110.100 162.600 110.200 ;
        RECT 157.400 109.800 162.600 110.100 ;
        RECT 6.200 109.100 6.600 109.200 ;
        RECT 12.600 109.100 13.000 109.200 ;
        RECT 16.600 109.100 17.000 109.200 ;
        RECT 24.600 109.100 25.000 109.200 ;
        RECT 30.200 109.100 30.600 109.200 ;
        RECT 6.200 108.800 30.600 109.100 ;
        RECT 39.000 109.100 39.400 109.200 ;
        RECT 46.200 109.100 46.600 109.200 ;
        RECT 39.000 108.800 46.600 109.100 ;
        RECT 109.400 109.100 109.800 109.200 ;
        RECT 110.200 109.100 110.600 109.200 ;
        RECT 109.400 108.800 110.600 109.100 ;
        RECT 162.200 109.100 162.600 109.200 ;
        RECT 168.600 109.100 169.000 109.200 ;
        RECT 162.200 108.800 169.000 109.100 ;
        RECT 20.600 108.100 21.000 108.200 ;
        RECT 27.800 108.100 28.200 108.200 ;
        RECT 20.600 107.800 28.200 108.100 ;
        RECT 43.000 108.100 43.400 108.200 ;
        RECT 55.000 108.100 55.400 108.200 ;
        RECT 43.000 107.800 55.400 108.100 ;
        RECT 55.800 108.100 56.200 108.200 ;
        RECT 57.400 108.100 57.800 108.200 ;
        RECT 97.400 108.100 97.800 108.200 ;
        RECT 55.800 107.800 57.800 108.100 ;
        RECT 58.200 107.800 97.800 108.100 ;
        RECT 134.200 108.100 134.600 108.200 ;
        RECT 143.800 108.100 144.200 108.200 ;
        RECT 134.200 107.800 144.200 108.100 ;
        RECT 166.200 107.800 166.600 108.200 ;
        RECT 11.800 107.100 12.200 107.200 ;
        RECT 13.400 107.100 13.800 107.200 ;
        RECT 19.800 107.100 20.200 107.200 ;
        RECT 11.800 106.800 20.200 107.100 ;
        RECT 41.400 107.100 41.800 107.200 ;
        RECT 42.200 107.100 42.600 107.200 ;
        RECT 41.400 106.800 42.600 107.100 ;
        RECT 46.200 107.100 46.600 107.200 ;
        RECT 52.600 107.100 53.000 107.200 ;
        RECT 46.200 106.800 53.000 107.100 ;
        RECT 57.400 107.100 57.800 107.200 ;
        RECT 58.200 107.100 58.500 107.800 ;
        RECT 166.200 107.200 166.500 107.800 ;
        RECT 57.400 106.800 58.500 107.100 ;
        RECT 77.400 107.100 77.800 107.200 ;
        RECT 78.200 107.100 78.600 107.200 ;
        RECT 77.400 106.800 78.600 107.100 ;
        RECT 82.200 107.100 82.600 107.200 ;
        RECT 83.800 107.100 84.200 107.200 ;
        RECT 82.200 106.800 84.200 107.100 ;
        RECT 86.200 107.100 86.600 107.200 ;
        RECT 107.000 107.100 107.400 107.200 ;
        RECT 86.200 106.800 107.400 107.100 ;
        RECT 126.200 107.100 126.600 107.200 ;
        RECT 143.000 107.100 143.400 107.200 ;
        RECT 146.200 107.100 146.600 107.200 ;
        RECT 147.000 107.100 147.400 107.200 ;
        RECT 126.200 106.800 131.300 107.100 ;
        RECT 143.000 106.800 147.400 107.100 ;
        RECT 147.800 107.100 148.200 107.200 ;
        RECT 149.400 107.100 149.800 107.200 ;
        RECT 147.800 106.800 149.800 107.100 ;
        RECT 163.000 107.100 163.400 107.200 ;
        RECT 163.800 107.100 164.200 107.200 ;
        RECT 163.000 106.800 164.200 107.100 ;
        RECT 164.600 106.800 165.000 107.200 ;
        RECT 166.200 106.800 166.600 107.200 ;
        RECT 168.600 107.100 169.000 107.200 ;
        RECT 170.200 107.100 170.600 107.200 ;
        RECT 168.600 106.800 170.600 107.100 ;
        RECT 131.000 106.200 131.300 106.800 ;
        RECT 12.600 106.100 13.000 106.200 ;
        RECT 3.800 105.800 13.000 106.100 ;
        RECT 22.200 106.100 22.600 106.200 ;
        RECT 42.200 106.100 42.600 106.200 ;
        RECT 61.400 106.100 61.800 106.200 ;
        RECT 22.200 105.800 61.800 106.100 ;
        RECT 63.800 106.100 64.200 106.200 ;
        RECT 65.400 106.100 65.800 106.200 ;
        RECT 63.800 105.800 65.800 106.100 ;
        RECT 99.000 106.100 99.400 106.200 ;
        RECT 99.800 106.100 100.200 106.200 ;
        RECT 103.000 106.100 103.400 106.200 ;
        RECT 99.000 105.800 103.400 106.100 ;
        RECT 112.600 106.100 113.000 106.200 ;
        RECT 115.800 106.100 116.200 106.200 ;
        RECT 112.600 105.800 116.200 106.100 ;
        RECT 131.000 105.800 131.400 106.200 ;
        RECT 143.800 105.800 144.200 106.200 ;
        RECT 148.600 106.100 149.000 106.200 ;
        RECT 155.000 106.100 155.400 106.200 ;
        RECT 161.400 106.100 161.800 106.200 ;
        RECT 162.200 106.100 162.600 106.200 ;
        RECT 148.600 105.800 160.100 106.100 ;
        RECT 161.400 105.800 162.600 106.100 ;
        RECT 164.600 106.100 164.900 106.800 ;
        RECT 167.800 106.100 168.200 106.200 ;
        RECT 169.400 106.100 169.800 106.200 ;
        RECT 164.600 105.800 169.800 106.100 ;
        RECT 173.400 106.100 173.800 106.200 ;
        RECT 175.800 106.100 176.200 106.200 ;
        RECT 173.400 105.800 176.200 106.100 ;
        RECT 3.800 105.200 4.100 105.800 ;
        RECT 143.800 105.200 144.100 105.800 ;
        RECT 159.800 105.200 160.100 105.800 ;
        RECT 3.800 104.800 4.200 105.200 ;
        RECT 32.600 105.100 33.000 105.200 ;
        RECT 47.800 105.100 48.200 105.200 ;
        RECT 51.000 105.100 51.400 105.200 ;
        RECT 32.600 104.800 43.300 105.100 ;
        RECT 47.800 104.800 51.400 105.100 ;
        RECT 55.800 105.100 56.200 105.200 ;
        RECT 56.600 105.100 57.000 105.200 ;
        RECT 60.600 105.100 61.000 105.200 ;
        RECT 55.800 104.800 61.000 105.100 ;
        RECT 63.800 105.100 64.200 105.200 ;
        RECT 64.600 105.100 65.000 105.200 ;
        RECT 63.800 104.800 65.000 105.100 ;
        RECT 143.800 104.800 144.200 105.200 ;
        RECT 159.800 104.800 160.200 105.200 ;
        RECT 165.400 105.100 165.800 105.200 ;
        RECT 167.000 105.100 167.400 105.200 ;
        RECT 165.400 104.800 167.400 105.100 ;
        RECT 43.000 104.200 43.300 104.800 ;
        RECT 27.800 103.800 28.200 104.200 ;
        RECT 40.600 104.100 41.000 104.200 ;
        RECT 41.400 104.100 41.800 104.200 ;
        RECT 40.600 103.800 41.800 104.100 ;
        RECT 43.000 103.800 43.400 104.200 ;
        RECT 51.000 104.100 51.400 104.200 ;
        RECT 45.400 103.800 51.400 104.100 ;
        RECT 64.600 104.100 65.000 104.200 ;
        RECT 100.600 104.100 101.000 104.200 ;
        RECT 64.600 103.800 101.000 104.100 ;
        RECT 120.600 104.100 121.000 104.200 ;
        RECT 123.000 104.100 123.400 104.200 ;
        RECT 120.600 103.800 123.400 104.100 ;
        RECT 9.400 102.800 9.800 103.200 ;
        RECT 27.800 103.100 28.100 103.800 ;
        RECT 45.400 103.100 45.700 103.800 ;
        RECT 27.800 102.800 45.700 103.100 ;
        RECT 46.200 103.100 46.600 103.200 ;
        RECT 48.600 103.100 49.000 103.200 ;
        RECT 46.200 102.800 49.000 103.100 ;
        RECT 49.400 103.100 49.800 103.200 ;
        RECT 51.000 103.100 51.400 103.200 ;
        RECT 49.400 102.800 51.400 103.100 ;
        RECT 63.000 102.800 63.400 103.200 ;
        RECT 79.000 103.100 79.400 103.200 ;
        RECT 135.000 103.100 135.400 103.200 ;
        RECT 79.000 102.800 135.400 103.100 ;
        RECT 9.400 102.100 9.700 102.800 ;
        RECT 15.000 102.100 15.400 102.200 ;
        RECT 9.400 101.800 15.400 102.100 ;
        RECT 32.600 102.100 33.000 102.200 ;
        RECT 63.000 102.100 63.300 102.800 ;
        RECT 32.600 101.800 63.300 102.100 ;
        RECT 67.800 102.100 68.200 102.200 ;
        RECT 83.000 102.100 83.400 102.200 ;
        RECT 67.800 101.800 83.400 102.100 ;
        RECT 85.400 102.100 85.800 102.200 ;
        RECT 96.600 102.100 97.000 102.200 ;
        RECT 113.400 102.100 113.800 102.200 ;
        RECT 85.400 101.800 113.800 102.100 ;
        RECT 128.600 102.100 129.000 102.200 ;
        RECT 129.400 102.100 129.800 102.200 ;
        RECT 128.600 101.800 129.800 102.100 ;
        RECT 163.000 102.100 163.400 102.200 ;
        RECT 165.400 102.100 165.800 102.200 ;
        RECT 163.000 101.800 165.800 102.100 ;
        RECT 42.200 101.100 42.600 101.200 ;
        RECT 47.800 101.100 48.200 101.200 ;
        RECT 42.200 100.800 48.200 101.100 ;
        RECT 61.400 101.100 61.800 101.200 ;
        RECT 76.600 101.100 77.000 101.200 ;
        RECT 98.200 101.100 98.600 101.200 ;
        RECT 133.400 101.100 133.800 101.200 ;
        RECT 61.400 100.800 133.800 101.100 ;
        RECT 147.000 101.100 147.400 101.200 ;
        RECT 163.000 101.100 163.400 101.200 ;
        RECT 147.000 100.800 163.400 101.100 ;
        RECT 45.400 100.100 45.800 100.200 ;
        RECT 73.400 100.100 73.800 100.200 ;
        RECT 45.400 99.800 73.800 100.100 ;
        RECT 86.200 99.800 86.600 100.200 ;
        RECT 153.400 100.100 153.800 100.200 ;
        RECT 159.000 100.100 159.400 100.200 ;
        RECT 153.400 99.800 159.400 100.100 ;
        RECT 86.200 99.200 86.500 99.800 ;
        RECT 15.800 99.100 16.200 99.200 ;
        RECT 42.200 99.100 42.600 99.200 ;
        RECT 15.800 98.800 42.600 99.100 ;
        RECT 86.200 98.800 86.600 99.200 ;
        RECT 91.000 99.100 91.400 99.200 ;
        RECT 94.200 99.100 94.600 99.200 ;
        RECT 99.800 99.100 100.200 99.200 ;
        RECT 91.000 98.800 100.200 99.100 ;
        RECT 114.200 98.800 114.600 99.200 ;
        RECT 133.400 99.100 133.800 99.200 ;
        RECT 159.800 99.100 160.200 99.200 ;
        RECT 164.600 99.100 165.000 99.200 ;
        RECT 133.400 98.800 165.000 99.100 ;
        RECT 114.200 98.200 114.500 98.800 ;
        RECT 9.400 97.800 9.800 98.200 ;
        RECT 13.400 98.100 13.800 98.200 ;
        RECT 18.200 98.100 18.600 98.200 ;
        RECT 13.400 97.800 18.600 98.100 ;
        RECT 19.000 98.100 19.400 98.200 ;
        RECT 19.800 98.100 20.200 98.200 ;
        RECT 40.600 98.100 41.000 98.200 ;
        RECT 19.000 97.800 41.000 98.100 ;
        RECT 45.400 98.100 45.800 98.200 ;
        RECT 46.200 98.100 46.600 98.200 ;
        RECT 45.400 97.800 46.600 98.100 ;
        RECT 50.200 98.100 50.600 98.200 ;
        RECT 87.800 98.100 88.200 98.200 ;
        RECT 50.200 97.800 88.200 98.100 ;
        RECT 114.200 97.800 114.600 98.200 ;
        RECT 9.400 97.100 9.700 97.800 ;
        RECT 35.800 97.100 36.200 97.200 ;
        RECT 9.400 96.800 36.200 97.100 ;
        RECT 38.200 97.100 38.600 97.200 ;
        RECT 39.800 97.100 40.200 97.200 ;
        RECT 48.600 97.100 49.000 97.200 ;
        RECT 38.200 96.800 49.000 97.100 ;
        RECT 55.800 97.100 56.200 97.200 ;
        RECT 62.200 97.100 62.600 97.200 ;
        RECT 55.800 96.800 62.600 97.100 ;
        RECT 64.600 97.100 65.000 97.200 ;
        RECT 76.600 97.100 77.000 97.200 ;
        RECT 64.600 96.800 77.000 97.100 ;
        RECT 81.400 97.100 81.800 97.200 ;
        RECT 99.800 97.100 100.200 97.200 ;
        RECT 104.600 97.100 105.000 97.200 ;
        RECT 81.400 96.800 105.000 97.100 ;
        RECT 160.600 96.800 161.000 97.200 ;
        RECT 15.000 96.100 15.400 96.200 ;
        RECT 16.600 96.100 17.000 96.200 ;
        RECT 15.000 95.800 17.000 96.100 ;
        RECT 23.800 96.100 24.200 96.200 ;
        RECT 30.200 96.100 30.600 96.200 ;
        RECT 23.800 95.800 30.600 96.100 ;
        RECT 33.400 96.100 33.800 96.200 ;
        RECT 36.600 96.100 37.000 96.200 ;
        RECT 47.000 96.100 47.400 96.200 ;
        RECT 47.800 96.100 48.200 96.200 ;
        RECT 33.400 95.800 48.200 96.100 ;
        RECT 73.400 95.800 73.800 96.200 ;
        RECT 91.800 96.100 92.200 96.200 ;
        RECT 95.800 96.100 96.200 96.200 ;
        RECT 96.600 96.100 97.000 96.200 ;
        RECT 91.800 95.800 97.000 96.100 ;
        RECT 160.600 96.100 160.900 96.800 ;
        RECT 171.000 96.100 171.400 96.200 ;
        RECT 160.600 95.800 171.400 96.100 ;
        RECT 3.000 95.100 3.400 95.200 ;
        RECT 11.800 95.100 12.200 95.200 ;
        RECT 3.000 94.800 12.200 95.100 ;
        RECT 12.600 95.100 13.000 95.200 ;
        RECT 14.200 95.100 14.600 95.200 ;
        RECT 12.600 94.800 14.600 95.100 ;
        RECT 21.400 95.100 21.800 95.200 ;
        RECT 24.600 95.100 25.000 95.200 ;
        RECT 21.400 94.800 25.000 95.100 ;
        RECT 29.400 95.100 29.800 95.200 ;
        RECT 42.200 95.100 42.600 95.200 ;
        RECT 47.000 95.100 47.400 95.200 ;
        RECT 59.800 95.100 60.200 95.200 ;
        RECT 29.400 94.800 60.200 95.100 ;
        RECT 63.000 95.100 63.400 95.200 ;
        RECT 70.200 95.100 70.600 95.200 ;
        RECT 63.000 94.800 70.600 95.100 ;
        RECT 73.400 95.100 73.700 95.800 ;
        RECT 91.800 95.100 92.200 95.200 ;
        RECT 73.400 94.800 92.200 95.100 ;
        RECT 100.600 95.100 101.000 95.200 ;
        RECT 106.200 95.100 106.600 95.200 ;
        RECT 100.600 94.800 106.600 95.100 ;
        RECT 107.000 95.100 107.400 95.200 ;
        RECT 112.600 95.100 113.000 95.200 ;
        RECT 113.400 95.100 113.800 95.200 ;
        RECT 107.000 94.800 113.800 95.100 ;
        RECT 122.200 95.100 122.600 95.200 ;
        RECT 159.000 95.100 159.400 95.200 ;
        RECT 163.800 95.100 164.200 95.200 ;
        RECT 122.200 94.800 159.400 95.100 ;
        RECT 162.200 94.800 164.200 95.100 ;
        RECT 158.200 94.200 158.500 94.800 ;
        RECT 162.200 94.200 162.500 94.800 ;
        RECT 10.200 94.100 10.600 94.200 ;
        RECT 19.800 94.100 20.200 94.200 ;
        RECT 25.400 94.100 25.800 94.200 ;
        RECT 10.200 93.800 25.800 94.100 ;
        RECT 42.200 94.100 42.600 94.200 ;
        RECT 44.600 94.100 45.000 94.200 ;
        RECT 42.200 93.800 45.000 94.100 ;
        RECT 45.400 94.100 45.800 94.200 ;
        RECT 46.200 94.100 46.600 94.200 ;
        RECT 45.400 93.800 46.600 94.100 ;
        RECT 53.400 94.100 53.800 94.200 ;
        RECT 55.800 94.100 56.200 94.200 ;
        RECT 53.400 93.800 56.200 94.100 ;
        RECT 73.400 94.100 73.800 94.200 ;
        RECT 80.600 94.100 81.000 94.200 ;
        RECT 92.600 94.100 93.000 94.200 ;
        RECT 73.400 93.800 81.000 94.100 ;
        RECT 83.000 93.800 93.000 94.100 ;
        RECT 96.600 94.100 97.000 94.200 ;
        RECT 104.600 94.100 105.000 94.200 ;
        RECT 96.600 93.800 105.000 94.100 ;
        RECT 112.600 94.100 113.000 94.200 ;
        RECT 115.000 94.100 115.400 94.200 ;
        RECT 137.400 94.100 137.800 94.200 ;
        RECT 112.600 93.800 137.800 94.100 ;
        RECT 158.200 93.800 158.600 94.200 ;
        RECT 162.200 93.800 162.600 94.200 ;
        RECT 83.000 93.200 83.300 93.800 ;
        RECT 20.600 93.100 21.000 93.200 ;
        RECT 24.600 93.100 25.000 93.200 ;
        RECT 31.800 93.100 32.200 93.200 ;
        RECT 43.000 93.100 43.400 93.200 ;
        RECT 20.600 92.800 22.500 93.100 ;
        RECT 24.600 92.800 43.400 93.100 ;
        RECT 45.400 93.100 45.800 93.200 ;
        RECT 55.800 93.100 56.200 93.200 ;
        RECT 45.400 92.800 56.200 93.100 ;
        RECT 57.400 93.100 57.800 93.200 ;
        RECT 58.200 93.100 58.600 93.200 ;
        RECT 57.400 92.800 58.600 93.100 ;
        RECT 83.000 92.800 83.400 93.200 ;
        RECT 95.800 93.100 96.200 93.200 ;
        RECT 98.200 93.100 98.600 93.200 ;
        RECT 95.800 92.800 98.600 93.100 ;
        RECT 117.400 93.100 117.800 93.200 ;
        RECT 175.000 93.100 175.400 93.200 ;
        RECT 117.400 92.800 175.400 93.100 ;
        RECT 22.200 92.200 22.500 92.800 ;
        RECT 22.200 92.100 22.600 92.200 ;
        RECT 25.400 92.100 25.800 92.200 ;
        RECT 22.200 91.800 25.800 92.100 ;
        RECT 40.600 92.100 41.000 92.200 ;
        RECT 42.200 92.100 42.600 92.200 ;
        RECT 46.200 92.100 46.600 92.200 ;
        RECT 40.600 91.800 46.600 92.100 ;
        RECT 55.000 92.100 55.400 92.200 ;
        RECT 59.800 92.100 60.200 92.200 ;
        RECT 55.000 91.800 60.200 92.100 ;
        RECT 74.200 92.100 74.600 92.200 ;
        RECT 75.800 92.100 76.200 92.200 ;
        RECT 99.800 92.100 100.200 92.200 ;
        RECT 74.200 91.800 100.200 92.100 ;
        RECT 115.800 92.100 116.200 92.200 ;
        RECT 127.800 92.100 128.200 92.200 ;
        RECT 115.800 91.800 128.200 92.100 ;
        RECT 135.800 92.100 136.200 92.200 ;
        RECT 143.000 92.100 143.400 92.200 ;
        RECT 135.800 91.800 143.400 92.100 ;
        RECT 147.000 92.100 147.400 92.200 ;
        RECT 164.600 92.100 165.000 92.200 ;
        RECT 147.000 91.800 165.000 92.100 ;
        RECT 166.200 92.100 166.600 92.200 ;
        RECT 173.400 92.100 173.800 92.200 ;
        RECT 166.200 91.800 173.800 92.100 ;
        RECT 37.400 91.100 37.800 91.200 ;
        RECT 64.600 91.100 65.000 91.200 ;
        RECT 37.400 90.800 65.000 91.100 ;
        RECT 123.800 91.100 124.200 91.200 ;
        RECT 129.400 91.100 129.800 91.200 ;
        RECT 123.800 90.800 129.800 91.100 ;
        RECT 140.600 91.100 141.000 91.200 ;
        RECT 152.600 91.100 153.000 91.200 ;
        RECT 177.400 91.100 177.800 91.200 ;
        RECT 140.600 90.800 177.800 91.100 ;
        RECT 11.800 90.100 12.200 90.200 ;
        RECT 21.400 90.100 21.800 90.200 ;
        RECT 11.800 89.800 21.800 90.100 ;
        RECT 51.800 90.100 52.200 90.200 ;
        RECT 59.800 90.100 60.200 90.200 ;
        RECT 51.800 89.800 60.200 90.100 ;
        RECT 70.200 90.100 70.600 90.200 ;
        RECT 75.000 90.100 75.400 90.200 ;
        RECT 70.200 89.800 75.400 90.100 ;
        RECT 99.800 90.100 100.200 90.200 ;
        RECT 102.200 90.100 102.600 90.200 ;
        RECT 99.800 89.800 102.600 90.100 ;
        RECT 150.200 90.100 150.600 90.200 ;
        RECT 151.000 90.100 151.400 90.200 ;
        RECT 150.200 89.800 151.400 90.100 ;
        RECT 10.200 89.100 10.600 89.200 ;
        RECT 15.000 89.100 15.400 89.200 ;
        RECT 10.200 88.800 15.400 89.100 ;
        RECT 25.400 89.100 25.800 89.200 ;
        RECT 28.600 89.100 29.000 89.200 ;
        RECT 25.400 88.800 29.000 89.100 ;
        RECT 47.800 89.100 48.200 89.200 ;
        RECT 51.800 89.100 52.200 89.200 ;
        RECT 47.800 88.800 52.200 89.100 ;
        RECT 53.400 89.100 53.800 89.200 ;
        RECT 59.000 89.100 59.400 89.200 ;
        RECT 53.400 88.800 59.400 89.100 ;
        RECT 59.800 89.100 60.200 89.200 ;
        RECT 62.200 89.100 62.600 89.200 ;
        RECT 83.000 89.100 83.400 89.200 ;
        RECT 59.800 88.800 83.400 89.100 ;
        RECT 83.800 89.100 84.200 89.200 ;
        RECT 115.000 89.100 115.400 89.200 ;
        RECT 83.800 88.800 115.400 89.100 ;
        RECT 147.800 89.100 148.200 89.200 ;
        RECT 161.400 89.100 161.800 89.200 ;
        RECT 147.800 88.800 161.800 89.100 ;
        RECT 163.000 89.100 163.400 89.200 ;
        RECT 163.800 89.100 164.200 89.200 ;
        RECT 163.000 88.800 164.200 89.100 ;
        RECT 167.000 88.800 167.400 89.200 ;
        RECT 11.000 88.100 11.400 88.200 ;
        RECT 14.200 88.100 14.600 88.200 ;
        RECT 11.000 87.800 14.600 88.100 ;
        RECT 17.400 88.100 17.800 88.200 ;
        RECT 20.600 88.100 21.000 88.200 ;
        RECT 27.000 88.100 27.400 88.200 ;
        RECT 56.600 88.100 57.000 88.200 ;
        RECT 67.800 88.100 68.200 88.200 ;
        RECT 17.400 87.800 43.300 88.100 ;
        RECT 56.600 87.800 68.200 88.100 ;
        RECT 69.400 88.100 69.800 88.200 ;
        RECT 93.400 88.100 93.800 88.200 ;
        RECT 102.200 88.100 102.600 88.200 ;
        RECT 69.400 87.800 93.800 88.100 ;
        RECT 94.200 87.800 102.600 88.100 ;
        RECT 144.600 88.100 145.000 88.200 ;
        RECT 158.200 88.100 158.600 88.200 ;
        RECT 163.800 88.100 164.200 88.200 ;
        RECT 144.600 87.800 149.700 88.100 ;
        RECT 158.200 87.800 164.200 88.100 ;
        RECT 167.000 88.100 167.300 88.800 ;
        RECT 171.000 88.100 171.400 88.200 ;
        RECT 167.000 87.800 171.400 88.100 ;
        RECT 172.600 88.100 173.000 88.200 ;
        RECT 173.400 88.100 173.800 88.200 ;
        RECT 172.600 87.800 173.800 88.100 ;
        RECT 174.200 88.100 174.600 88.200 ;
        RECT 179.800 88.100 180.200 88.200 ;
        RECT 174.200 87.800 180.200 88.100 ;
        RECT 43.000 87.200 43.300 87.800 ;
        RECT 19.800 87.100 20.200 87.200 ;
        RECT 22.200 87.100 22.600 87.200 ;
        RECT 29.400 87.100 29.800 87.200 ;
        RECT 19.800 86.800 29.800 87.100 ;
        RECT 43.000 87.100 43.400 87.200 ;
        RECT 43.800 87.100 44.200 87.200 ;
        RECT 43.000 86.800 44.200 87.100 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 56.600 86.800 57.000 87.200 ;
        RECT 66.200 87.100 66.600 87.200 ;
        RECT 68.600 87.100 69.000 87.200 ;
        RECT 66.200 86.800 69.000 87.100 ;
        RECT 77.400 86.800 77.800 87.200 ;
        RECT 84.600 87.100 85.000 87.200 ;
        RECT 94.200 87.100 94.500 87.800 ;
        RECT 149.400 87.200 149.700 87.800 ;
        RECT 84.600 86.800 94.500 87.100 ;
        RECT 95.000 87.100 95.400 87.200 ;
        RECT 99.000 87.100 99.400 87.200 ;
        RECT 95.000 86.800 99.400 87.100 ;
        RECT 101.400 87.100 101.800 87.200 ;
        RECT 106.200 87.100 106.600 87.200 ;
        RECT 101.400 86.800 106.600 87.100 ;
        RECT 116.600 86.800 117.000 87.200 ;
        RECT 149.400 86.800 149.800 87.200 ;
        RECT 159.000 87.100 159.400 87.200 ;
        RECT 159.800 87.100 160.200 87.200 ;
        RECT 159.000 86.800 160.200 87.100 ;
        RECT 163.800 87.100 164.200 87.200 ;
        RECT 178.200 87.100 178.600 87.200 ;
        RECT 163.800 86.800 178.600 87.100 ;
        RECT 44.600 86.200 44.900 86.800 ;
        RECT 3.000 86.100 3.400 86.200 ;
        RECT 10.200 86.100 10.600 86.200 ;
        RECT 3.000 85.800 10.600 86.100 ;
        RECT 17.400 86.100 17.800 86.200 ;
        RECT 23.800 86.100 24.200 86.200 ;
        RECT 17.400 85.800 24.200 86.100 ;
        RECT 25.400 86.100 25.800 86.200 ;
        RECT 26.200 86.100 26.600 86.200 ;
        RECT 25.400 85.800 26.600 86.100 ;
        RECT 33.400 86.100 33.800 86.200 ;
        RECT 34.200 86.100 34.600 86.200 ;
        RECT 33.400 85.800 34.600 86.100 ;
        RECT 35.000 86.100 35.400 86.200 ;
        RECT 43.800 86.100 44.200 86.200 ;
        RECT 35.000 85.800 44.200 86.100 ;
        RECT 44.600 85.800 45.000 86.200 ;
        RECT 47.800 86.100 48.200 86.200 ;
        RECT 56.600 86.100 56.900 86.800 ;
        RECT 77.400 86.200 77.700 86.800 ;
        RECT 116.600 86.200 116.900 86.800 ;
        RECT 47.800 85.800 56.900 86.100 ;
        RECT 57.400 86.100 57.800 86.200 ;
        RECT 62.200 86.100 62.600 86.200 ;
        RECT 67.800 86.100 68.200 86.200 ;
        RECT 70.200 86.100 70.600 86.200 ;
        RECT 57.400 85.800 65.700 86.100 ;
        RECT 67.800 85.800 70.600 86.100 ;
        RECT 77.400 85.800 77.800 86.200 ;
        RECT 83.000 86.100 83.400 86.200 ;
        RECT 95.800 86.100 96.200 86.200 ;
        RECT 83.000 85.800 96.200 86.100 ;
        RECT 97.400 86.100 97.800 86.200 ;
        RECT 98.200 86.100 98.600 86.200 ;
        RECT 97.400 85.800 98.600 86.100 ;
        RECT 99.000 86.100 99.400 86.200 ;
        RECT 103.000 86.100 103.400 86.200 ;
        RECT 99.000 85.800 103.400 86.100 ;
        RECT 116.600 85.800 117.000 86.200 ;
        RECT 123.000 86.100 123.400 86.200 ;
        RECT 125.400 86.100 125.800 86.200 ;
        RECT 123.000 85.800 125.800 86.100 ;
        RECT 166.200 86.100 166.600 86.200 ;
        RECT 168.600 86.100 169.000 86.200 ;
        RECT 166.200 85.800 169.000 86.100 ;
        RECT 170.200 86.100 170.600 86.200 ;
        RECT 171.000 86.100 171.400 86.200 ;
        RECT 170.200 85.800 171.400 86.100 ;
        RECT 18.200 85.100 18.600 85.200 ;
        RECT 19.000 85.100 19.400 85.200 ;
        RECT 18.200 84.800 19.400 85.100 ;
        RECT 27.800 85.100 28.200 85.200 ;
        RECT 40.600 85.100 41.000 85.200 ;
        RECT 52.600 85.100 53.000 85.200 ;
        RECT 27.800 84.800 53.000 85.100 ;
        RECT 63.800 85.100 64.200 85.200 ;
        RECT 64.600 85.100 65.000 85.200 ;
        RECT 63.800 84.800 65.000 85.100 ;
        RECT 65.400 85.100 65.700 85.800 ;
        RECT 95.000 85.100 95.400 85.200 ;
        RECT 65.400 84.800 95.400 85.100 ;
        RECT 115.800 85.100 116.200 85.200 ;
        RECT 117.400 85.100 117.800 85.200 ;
        RECT 115.800 84.800 117.800 85.100 ;
        RECT 119.000 85.100 119.400 85.200 ;
        RECT 123.000 85.100 123.400 85.200 ;
        RECT 119.000 84.800 123.400 85.100 ;
        RECT 137.400 85.100 137.800 85.200 ;
        RECT 155.000 85.100 155.400 85.200 ;
        RECT 162.200 85.100 162.600 85.200 ;
        RECT 170.200 85.100 170.600 85.200 ;
        RECT 171.800 85.100 172.200 85.200 ;
        RECT 137.400 84.800 172.200 85.100 ;
        RECT 46.200 84.200 46.500 84.800 ;
        RECT 21.400 84.100 21.800 84.200 ;
        RECT 23.800 84.100 24.200 84.200 ;
        RECT 21.400 83.800 24.200 84.100 ;
        RECT 25.400 84.100 25.800 84.200 ;
        RECT 30.200 84.100 30.600 84.200 ;
        RECT 25.400 83.800 30.600 84.100 ;
        RECT 35.000 84.100 35.400 84.200 ;
        RECT 39.000 84.100 39.400 84.200 ;
        RECT 35.000 83.800 39.400 84.100 ;
        RECT 44.600 84.100 45.000 84.200 ;
        RECT 45.400 84.100 45.800 84.200 ;
        RECT 44.600 83.800 45.800 84.100 ;
        RECT 46.200 83.800 46.600 84.200 ;
        RECT 64.600 84.100 65.000 84.200 ;
        RECT 69.400 84.100 69.800 84.200 ;
        RECT 76.600 84.100 77.000 84.200 ;
        RECT 64.600 83.800 77.000 84.100 ;
        RECT 80.600 84.100 81.000 84.200 ;
        RECT 87.000 84.100 87.400 84.200 ;
        RECT 80.600 83.800 87.400 84.100 ;
        RECT 93.400 84.100 93.800 84.200 ;
        RECT 96.600 84.100 97.000 84.200 ;
        RECT 114.200 84.100 114.600 84.200 ;
        RECT 93.400 83.800 114.600 84.100 ;
        RECT 167.000 84.100 167.400 84.200 ;
        RECT 175.000 84.100 175.400 84.200 ;
        RECT 167.000 83.800 175.400 84.100 ;
        RECT 27.800 82.800 28.200 83.200 ;
        RECT 56.600 83.100 57.000 83.200 ;
        RECT 75.000 83.100 75.400 83.200 ;
        RECT 56.600 82.800 75.400 83.100 ;
        RECT 27.800 82.200 28.100 82.800 ;
        RECT 27.800 82.100 28.200 82.200 ;
        RECT 39.800 82.100 40.200 82.200 ;
        RECT 43.000 82.100 43.400 82.200 ;
        RECT 27.800 81.800 43.400 82.100 ;
        RECT 66.200 82.100 66.600 82.200 ;
        RECT 69.400 82.100 69.800 82.200 ;
        RECT 66.200 81.800 69.800 82.100 ;
        RECT 71.800 82.100 72.200 82.200 ;
        RECT 74.200 82.100 74.600 82.200 ;
        RECT 100.600 82.100 101.000 82.200 ;
        RECT 71.800 81.800 101.000 82.100 ;
        RECT 131.800 82.100 132.200 82.200 ;
        RECT 132.600 82.100 133.000 82.200 ;
        RECT 131.800 81.800 133.000 82.100 ;
        RECT 75.800 81.100 76.200 81.200 ;
        RECT 120.600 81.100 121.000 81.200 ;
        RECT 75.800 80.800 121.000 81.100 ;
        RECT 127.800 81.100 128.200 81.200 ;
        RECT 133.400 81.100 133.800 81.200 ;
        RECT 127.800 80.800 133.800 81.100 ;
        RECT 39.000 80.100 39.400 80.200 ;
        RECT 53.400 80.100 53.800 80.200 ;
        RECT 39.000 79.800 53.800 80.100 ;
        RECT 72.600 80.100 73.000 80.200 ;
        RECT 75.800 80.100 76.100 80.800 ;
        RECT 72.600 79.800 76.100 80.100 ;
        RECT 100.600 80.100 101.000 80.200 ;
        RECT 132.600 80.100 133.000 80.200 ;
        RECT 135.800 80.100 136.200 80.200 ;
        RECT 100.600 79.800 136.200 80.100 ;
        RECT 26.200 79.100 26.600 79.200 ;
        RECT 78.200 79.100 78.600 79.200 ;
        RECT 91.000 79.100 91.400 79.200 ;
        RECT 26.200 78.800 74.500 79.100 ;
        RECT 78.200 78.800 91.400 79.100 ;
        RECT 102.200 79.100 102.600 79.200 ;
        RECT 111.000 79.100 111.400 79.200 ;
        RECT 114.200 79.100 114.600 79.200 ;
        RECT 102.200 78.800 114.600 79.100 ;
        RECT 170.200 79.100 170.600 79.200 ;
        RECT 171.000 79.100 171.400 79.200 ;
        RECT 170.200 78.800 171.400 79.100 ;
        RECT 74.200 78.200 74.500 78.800 ;
        RECT 12.600 77.800 13.000 78.200 ;
        RECT 19.800 78.100 20.200 78.200 ;
        RECT 22.200 78.100 22.600 78.200 ;
        RECT 28.600 78.100 29.000 78.200 ;
        RECT 19.800 77.800 29.000 78.100 ;
        RECT 39.000 78.100 39.400 78.200 ;
        RECT 43.800 78.100 44.200 78.200 ;
        RECT 51.800 78.100 52.200 78.200 ;
        RECT 39.000 77.800 52.200 78.100 ;
        RECT 63.000 78.100 63.400 78.200 ;
        RECT 73.400 78.100 73.800 78.200 ;
        RECT 63.000 77.800 73.800 78.100 ;
        RECT 74.200 77.800 74.600 78.200 ;
        RECT 83.000 78.100 83.400 78.200 ;
        RECT 86.200 78.100 86.600 78.200 ;
        RECT 97.400 78.100 97.800 78.200 ;
        RECT 83.000 77.800 97.800 78.100 ;
        RECT 102.200 78.100 102.600 78.200 ;
        RECT 105.400 78.100 105.800 78.200 ;
        RECT 102.200 77.800 105.800 78.100 ;
        RECT 108.600 78.100 109.000 78.200 ;
        RECT 114.200 78.100 114.600 78.200 ;
        RECT 122.200 78.100 122.600 78.200 ;
        RECT 108.600 77.800 122.600 78.100 ;
        RECT 123.800 78.100 124.200 78.200 ;
        RECT 139.000 78.100 139.400 78.200 ;
        RECT 123.800 77.800 139.400 78.100 ;
        RECT 12.600 77.100 12.900 77.800 ;
        RECT 23.800 77.100 24.200 77.200 ;
        RECT 12.600 76.800 24.200 77.100 ;
        RECT 55.800 77.100 56.200 77.200 ;
        RECT 63.800 77.100 64.200 77.200 ;
        RECT 55.800 76.800 64.200 77.100 ;
        RECT 73.400 77.100 73.800 77.200 ;
        RECT 87.000 77.100 87.400 77.200 ;
        RECT 73.400 76.800 87.400 77.100 ;
        RECT 93.400 77.100 93.800 77.200 ;
        RECT 100.600 77.100 101.000 77.200 ;
        RECT 111.800 77.100 112.200 77.200 ;
        RECT 93.400 76.800 112.200 77.100 ;
        RECT 112.600 77.100 113.000 77.200 ;
        RECT 113.400 77.100 113.800 77.200 ;
        RECT 112.600 76.800 113.800 77.100 ;
        RECT 118.200 77.100 118.600 77.200 ;
        RECT 123.800 77.100 124.200 77.200 ;
        RECT 118.200 76.800 124.200 77.100 ;
        RECT 124.600 77.100 125.000 77.200 ;
        RECT 128.600 77.100 129.000 77.200 ;
        RECT 124.600 76.800 129.000 77.100 ;
        RECT 131.000 77.100 131.400 77.200 ;
        RECT 137.400 77.100 137.800 77.200 ;
        RECT 131.000 76.800 137.800 77.100 ;
        RECT 19.000 76.100 19.400 76.200 ;
        RECT 21.400 76.100 21.800 76.200 ;
        RECT 23.000 76.100 23.400 76.200 ;
        RECT 49.400 76.100 49.800 76.200 ;
        RECT 50.200 76.100 50.600 76.200 ;
        RECT 19.000 75.800 20.900 76.100 ;
        RECT 21.400 75.800 23.400 76.100 ;
        RECT 45.400 75.800 50.600 76.100 ;
        RECT 55.000 76.100 55.400 76.200 ;
        RECT 61.400 76.100 61.800 76.200 ;
        RECT 55.000 75.800 61.800 76.100 ;
        RECT 66.200 76.100 66.600 76.200 ;
        RECT 91.800 76.100 92.200 76.200 ;
        RECT 132.600 76.100 133.000 76.200 ;
        RECT 66.200 75.800 133.000 76.100 ;
        RECT 135.000 75.800 135.400 76.200 ;
        RECT 143.000 75.800 143.400 76.200 ;
        RECT 165.400 75.800 165.800 76.200 ;
        RECT 3.000 75.100 3.400 75.200 ;
        RECT 15.800 75.100 16.200 75.200 ;
        RECT 3.000 74.800 16.200 75.100 ;
        RECT 20.600 75.100 20.900 75.800 ;
        RECT 45.400 75.200 45.700 75.800 ;
        RECT 23.000 75.100 23.400 75.200 ;
        RECT 20.600 74.800 23.400 75.100 ;
        RECT 30.200 75.100 30.600 75.200 ;
        RECT 37.400 75.100 37.800 75.200 ;
        RECT 30.200 74.800 37.800 75.100 ;
        RECT 45.400 74.800 45.800 75.200 ;
        RECT 50.200 75.100 50.600 75.200 ;
        RECT 63.800 75.100 64.200 75.200 ;
        RECT 50.200 74.800 64.200 75.100 ;
        RECT 69.400 75.100 69.800 75.200 ;
        RECT 75.000 75.100 75.400 75.200 ;
        RECT 69.400 74.800 75.400 75.100 ;
        RECT 84.600 74.800 85.000 75.200 ;
        RECT 99.800 75.100 100.200 75.200 ;
        RECT 107.000 75.100 107.400 75.200 ;
        RECT 114.200 75.100 114.600 75.200 ;
        RECT 127.000 75.100 127.400 75.200 ;
        RECT 128.600 75.100 129.000 75.200 ;
        RECT 99.800 74.800 129.000 75.100 ;
        RECT 129.400 75.100 129.800 75.200 ;
        RECT 133.400 75.100 133.800 75.200 ;
        RECT 129.400 74.800 133.800 75.100 ;
        RECT 135.000 75.100 135.300 75.800 ;
        RECT 143.000 75.200 143.300 75.800 ;
        RECT 142.200 75.100 142.600 75.200 ;
        RECT 135.000 74.800 142.600 75.100 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 157.400 75.100 157.800 75.200 ;
        RECT 162.200 75.100 162.600 75.200 ;
        RECT 165.400 75.100 165.700 75.800 ;
        RECT 157.400 74.800 165.700 75.100 ;
        RECT 168.600 75.100 169.000 75.200 ;
        RECT 175.000 75.100 175.400 75.200 ;
        RECT 168.600 74.800 175.400 75.100 ;
        RECT 84.600 74.200 84.900 74.800 ;
        RECT 9.400 74.100 9.800 74.200 ;
        RECT 14.200 74.100 14.600 74.200 ;
        RECT 9.400 73.800 14.600 74.100 ;
        RECT 57.400 74.100 57.800 74.200 ;
        RECT 67.800 74.100 68.200 74.200 ;
        RECT 57.400 73.800 68.200 74.100 ;
        RECT 82.200 74.100 82.600 74.200 ;
        RECT 83.000 74.100 83.400 74.200 ;
        RECT 82.200 73.800 83.400 74.100 ;
        RECT 84.600 73.800 85.000 74.200 ;
        RECT 96.600 74.100 97.000 74.200 ;
        RECT 97.400 74.100 97.800 74.200 ;
        RECT 96.600 73.800 97.800 74.100 ;
        RECT 106.200 74.100 106.600 74.200 ;
        RECT 143.800 74.100 144.200 74.200 ;
        RECT 166.200 74.100 166.600 74.200 ;
        RECT 174.200 74.100 174.600 74.200 ;
        RECT 106.200 73.800 174.600 74.100 ;
        RECT 3.800 73.100 4.200 73.200 ;
        RECT 11.800 73.100 12.200 73.200 ;
        RECT 3.800 72.800 12.200 73.100 ;
        RECT 15.000 73.100 15.400 73.200 ;
        RECT 20.600 73.100 21.000 73.200 ;
        RECT 15.000 72.800 21.000 73.100 ;
        RECT 63.000 73.100 63.400 73.200 ;
        RECT 70.200 73.100 70.600 73.200 ;
        RECT 63.000 72.800 70.600 73.100 ;
        RECT 100.600 73.100 101.000 73.200 ;
        RECT 102.200 73.100 102.600 73.200 ;
        RECT 116.600 73.100 117.000 73.200 ;
        RECT 100.600 72.800 117.000 73.100 ;
        RECT 119.000 72.800 119.400 73.200 ;
        RECT 132.600 73.100 133.000 73.200 ;
        RECT 140.600 73.100 141.000 73.200 ;
        RECT 132.600 72.800 141.000 73.100 ;
        RECT 144.600 73.100 145.000 73.200 ;
        RECT 144.600 72.800 156.100 73.100 ;
        RECT 119.000 72.200 119.300 72.800 ;
        RECT 155.800 72.200 156.100 72.800 ;
        RECT 6.200 72.100 6.600 72.200 ;
        RECT 15.800 72.100 16.200 72.200 ;
        RECT 6.200 71.800 16.200 72.100 ;
        RECT 43.800 72.100 44.200 72.200 ;
        RECT 54.200 72.100 54.600 72.200 ;
        RECT 59.800 72.100 60.200 72.200 ;
        RECT 43.800 71.800 60.200 72.100 ;
        RECT 70.200 72.100 70.600 72.200 ;
        RECT 78.200 72.100 78.600 72.200 ;
        RECT 70.200 71.800 78.600 72.100 ;
        RECT 81.400 72.100 81.800 72.200 ;
        RECT 85.400 72.100 85.800 72.200 ;
        RECT 81.400 71.800 85.800 72.100 ;
        RECT 110.200 72.100 110.600 72.200 ;
        RECT 117.400 72.100 117.800 72.200 ;
        RECT 110.200 71.800 117.800 72.100 ;
        RECT 119.000 71.800 119.400 72.200 ;
        RECT 134.200 72.100 134.600 72.200 ;
        RECT 147.000 72.100 147.400 72.200 ;
        RECT 134.200 71.800 147.400 72.100 ;
        RECT 155.800 71.800 156.200 72.200 ;
        RECT 168.600 72.100 169.000 72.200 ;
        RECT 175.800 72.100 176.200 72.200 ;
        RECT 163.800 71.800 176.200 72.100 ;
        RECT 163.800 71.200 164.100 71.800 ;
        RECT 57.400 71.100 57.800 71.200 ;
        RECT 77.400 71.100 77.800 71.200 ;
        RECT 84.600 71.100 85.000 71.200 ;
        RECT 57.400 70.800 85.000 71.100 ;
        RECT 95.000 71.100 95.400 71.200 ;
        RECT 99.800 71.100 100.200 71.200 ;
        RECT 95.000 70.800 100.200 71.100 ;
        RECT 103.800 71.100 104.200 71.200 ;
        RECT 118.200 71.100 118.600 71.200 ;
        RECT 103.800 70.800 118.600 71.100 ;
        RECT 123.800 71.100 124.200 71.200 ;
        RECT 138.200 71.100 138.600 71.200 ;
        RECT 153.400 71.100 153.800 71.200 ;
        RECT 123.800 70.800 153.800 71.100 ;
        RECT 155.000 70.800 155.400 71.200 ;
        RECT 163.800 70.800 164.200 71.200 ;
        RECT 155.000 70.200 155.300 70.800 ;
        RECT 8.600 70.100 9.000 70.200 ;
        RECT 10.200 70.100 10.600 70.200 ;
        RECT 8.600 69.800 10.600 70.100 ;
        RECT 55.000 70.100 55.400 70.200 ;
        RECT 55.800 70.100 56.200 70.200 ;
        RECT 55.000 69.800 56.200 70.100 ;
        RECT 64.600 70.100 65.000 70.200 ;
        RECT 72.600 70.100 73.000 70.200 ;
        RECT 110.200 70.100 110.600 70.200 ;
        RECT 127.000 70.100 127.400 70.200 ;
        RECT 64.600 69.800 73.000 70.100 ;
        RECT 98.200 69.800 127.400 70.100 ;
        RECT 155.000 69.800 155.400 70.200 ;
        RECT 98.200 69.200 98.500 69.800 ;
        RECT 10.200 69.100 10.600 69.200 ;
        RECT 11.000 69.100 11.400 69.200 ;
        RECT 10.200 68.800 11.400 69.100 ;
        RECT 18.200 69.100 18.600 69.200 ;
        RECT 28.600 69.100 29.000 69.200 ;
        RECT 18.200 68.800 29.000 69.100 ;
        RECT 48.600 69.100 49.000 69.200 ;
        RECT 79.800 69.100 80.200 69.200 ;
        RECT 86.200 69.100 86.600 69.200 ;
        RECT 48.600 68.800 67.300 69.100 ;
        RECT 79.800 68.800 86.600 69.100 ;
        RECT 92.600 69.100 93.000 69.200 ;
        RECT 98.200 69.100 98.600 69.200 ;
        RECT 92.600 68.800 98.600 69.100 ;
        RECT 99.800 69.100 100.200 69.200 ;
        RECT 101.400 69.100 101.800 69.200 ;
        RECT 99.800 68.800 101.800 69.100 ;
        RECT 107.800 69.100 108.200 69.200 ;
        RECT 111.000 69.100 111.400 69.200 ;
        RECT 107.800 68.800 111.400 69.100 ;
        RECT 111.800 69.100 112.200 69.200 ;
        RECT 141.400 69.100 141.800 69.200 ;
        RECT 111.800 68.800 141.800 69.100 ;
        RECT 154.200 69.100 154.600 69.200 ;
        RECT 156.600 69.100 157.000 69.200 ;
        RECT 154.200 68.800 157.000 69.100 ;
        RECT 158.200 69.100 158.600 69.200 ;
        RECT 163.800 69.100 164.200 69.200 ;
        RECT 167.000 69.100 167.400 69.200 ;
        RECT 158.200 68.800 164.200 69.100 ;
        RECT 164.600 68.800 167.400 69.100 ;
        RECT 67.000 68.200 67.300 68.800 ;
        RECT 164.600 68.200 164.900 68.800 ;
        RECT 25.400 68.100 25.800 68.200 ;
        RECT 26.200 68.100 26.600 68.200 ;
        RECT 27.800 68.100 28.200 68.200 ;
        RECT 25.400 67.800 28.200 68.100 ;
        RECT 28.600 68.100 29.000 68.200 ;
        RECT 48.600 68.100 49.000 68.200 ;
        RECT 53.400 68.100 53.800 68.200 ;
        RECT 56.600 68.100 57.000 68.200 ;
        RECT 28.600 67.800 57.000 68.100 ;
        RECT 67.000 67.800 67.400 68.200 ;
        RECT 91.000 68.100 91.400 68.200 ;
        RECT 91.000 67.800 101.700 68.100 ;
        RECT 101.400 67.200 101.700 67.800 ;
        RECT 116.600 67.800 117.000 68.200 ;
        RECT 121.400 68.100 121.800 68.200 ;
        RECT 135.800 68.100 136.200 68.200 ;
        RECT 121.400 67.800 136.200 68.100 ;
        RECT 143.800 68.100 144.200 68.200 ;
        RECT 161.400 68.100 161.800 68.200 ;
        RECT 143.800 67.800 161.800 68.100 ;
        RECT 163.000 67.800 163.400 68.200 ;
        RECT 164.600 67.800 165.000 68.200 ;
        RECT 116.600 67.200 116.900 67.800 ;
        RECT 5.400 67.100 5.800 67.200 ;
        RECT 19.800 67.100 20.200 67.200 ;
        RECT 5.400 66.800 20.200 67.100 ;
        RECT 22.200 67.100 22.600 67.200 ;
        RECT 26.200 67.100 26.600 67.200 ;
        RECT 22.200 66.800 26.600 67.100 ;
        RECT 42.200 66.800 42.600 67.200 ;
        RECT 45.400 67.100 45.800 67.200 ;
        RECT 51.000 67.100 51.400 67.200 ;
        RECT 45.400 66.800 51.400 67.100 ;
        RECT 54.200 67.100 54.600 67.200 ;
        RECT 55.000 67.100 55.400 67.200 ;
        RECT 54.200 66.800 55.400 67.100 ;
        RECT 62.200 67.100 62.600 67.200 ;
        RECT 63.800 67.100 64.200 67.200 ;
        RECT 62.200 66.800 64.200 67.100 ;
        RECT 67.800 66.800 68.200 67.200 ;
        RECT 72.600 67.100 73.000 67.200 ;
        RECT 85.400 67.100 85.800 67.200 ;
        RECT 91.800 67.100 92.200 67.200 ;
        RECT 72.600 66.800 92.200 67.100 ;
        RECT 98.200 67.100 98.600 67.200 ;
        RECT 99.800 67.100 100.200 67.200 ;
        RECT 98.200 66.800 100.200 67.100 ;
        RECT 101.400 66.800 101.800 67.200 ;
        RECT 103.000 67.100 103.400 67.200 ;
        RECT 103.800 67.100 104.200 67.200 ;
        RECT 103.000 66.800 104.200 67.100 ;
        RECT 107.000 66.800 107.400 67.200 ;
        RECT 116.600 66.800 117.000 67.200 ;
        RECT 117.400 67.100 117.800 67.200 ;
        RECT 121.400 67.100 121.800 67.200 ;
        RECT 117.400 66.800 121.800 67.100 ;
        RECT 123.800 67.100 124.200 67.200 ;
        RECT 134.200 67.100 134.600 67.200 ;
        RECT 123.800 66.800 134.600 67.100 ;
        RECT 141.400 67.100 141.800 67.200 ;
        RECT 163.000 67.100 163.300 67.800 ;
        RECT 167.800 67.100 168.200 67.200 ;
        RECT 141.400 66.800 168.200 67.100 ;
        RECT 7.800 66.100 8.200 66.200 ;
        RECT 14.200 66.100 14.600 66.200 ;
        RECT 21.400 66.100 21.800 66.200 ;
        RECT 7.800 65.800 14.600 66.100 ;
        RECT 19.000 65.800 21.800 66.100 ;
        RECT 23.800 66.100 24.200 66.200 ;
        RECT 32.600 66.100 33.000 66.200 ;
        RECT 23.800 65.800 33.000 66.100 ;
        RECT 38.200 66.100 38.600 66.200 ;
        RECT 42.200 66.100 42.500 66.800 ;
        RECT 67.800 66.200 68.100 66.800 ;
        RECT 38.200 65.800 42.500 66.100 ;
        RECT 43.000 66.100 43.400 66.200 ;
        RECT 49.400 66.100 49.800 66.200 ;
        RECT 66.200 66.100 66.600 66.200 ;
        RECT 43.000 65.800 66.600 66.100 ;
        RECT 67.800 65.800 68.200 66.200 ;
        RECT 74.200 66.100 74.600 66.200 ;
        RECT 81.400 66.100 81.800 66.200 ;
        RECT 74.200 65.800 81.800 66.100 ;
        RECT 85.400 65.800 85.800 66.200 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 87.000 66.100 87.400 66.200 ;
        RECT 107.000 66.100 107.300 66.800 ;
        RECT 87.000 65.800 107.300 66.100 ;
        RECT 117.400 66.100 117.800 66.200 ;
        RECT 118.200 66.100 118.600 66.200 ;
        RECT 117.400 65.800 118.600 66.100 ;
        RECT 123.000 66.100 123.400 66.200 ;
        RECT 135.000 66.100 135.400 66.200 ;
        RECT 135.800 66.100 136.200 66.200 ;
        RECT 123.000 65.800 127.300 66.100 ;
        RECT 135.000 65.800 136.200 66.100 ;
        RECT 140.600 66.100 141.000 66.200 ;
        RECT 160.600 66.100 161.000 66.200 ;
        RECT 140.600 65.800 161.000 66.100 ;
        RECT 161.400 66.100 161.800 66.200 ;
        RECT 164.600 66.100 165.000 66.200 ;
        RECT 161.400 65.800 165.000 66.100 ;
        RECT 167.800 66.100 168.200 66.200 ;
        RECT 172.600 66.100 173.000 66.200 ;
        RECT 167.800 65.800 173.000 66.100 ;
        RECT 19.000 65.200 19.300 65.800 ;
        RECT 85.400 65.200 85.700 65.800 ;
        RECT 86.200 65.200 86.500 65.800 ;
        RECT 127.000 65.200 127.300 65.800 ;
        RECT 19.000 64.800 19.400 65.200 ;
        RECT 19.800 65.100 20.200 65.200 ;
        RECT 20.600 65.100 21.000 65.200 ;
        RECT 19.800 64.800 21.000 65.100 ;
        RECT 59.800 65.100 60.200 65.200 ;
        RECT 83.000 65.100 83.400 65.200 ;
        RECT 59.800 64.800 83.400 65.100 ;
        RECT 85.400 64.800 85.800 65.200 ;
        RECT 86.200 64.800 86.600 65.200 ;
        RECT 91.800 65.100 92.200 65.200 ;
        RECT 105.400 65.100 105.800 65.200 ;
        RECT 115.800 65.100 116.200 65.200 ;
        RECT 119.800 65.100 120.200 65.200 ;
        RECT 91.800 64.800 120.200 65.100 ;
        RECT 127.000 64.800 127.400 65.200 ;
        RECT 143.000 65.100 143.400 65.200 ;
        RECT 147.800 65.100 148.200 65.200 ;
        RECT 143.000 64.800 148.200 65.100 ;
        RECT 151.800 65.100 152.200 65.200 ;
        RECT 152.600 65.100 153.000 65.200 ;
        RECT 151.800 64.800 153.000 65.100 ;
        RECT 155.000 65.100 155.400 65.200 ;
        RECT 167.000 65.100 167.400 65.200 ;
        RECT 168.600 65.100 169.000 65.200 ;
        RECT 155.000 64.800 169.000 65.100 ;
        RECT 19.000 64.100 19.400 64.200 ;
        RECT 56.600 64.100 57.000 64.200 ;
        RECT 19.000 63.800 57.000 64.100 ;
        RECT 60.600 64.100 61.000 64.200 ;
        RECT 72.600 64.100 73.000 64.200 ;
        RECT 60.600 63.800 73.000 64.100 ;
        RECT 84.600 64.100 85.000 64.200 ;
        RECT 95.800 64.100 96.200 64.200 ;
        RECT 106.200 64.100 106.600 64.200 ;
        RECT 84.600 63.800 106.600 64.100 ;
        RECT 145.400 64.100 145.800 64.200 ;
        RECT 146.200 64.100 146.600 64.200 ;
        RECT 145.400 63.800 146.600 64.100 ;
        RECT 159.800 64.100 160.200 64.200 ;
        RECT 163.000 64.100 163.400 64.200 ;
        RECT 159.800 63.800 163.400 64.100 ;
        RECT 43.000 63.100 43.400 63.200 ;
        RECT 43.800 63.100 44.200 63.200 ;
        RECT 43.000 62.800 44.200 63.100 ;
        RECT 47.800 63.100 48.200 63.200 ;
        RECT 78.200 63.100 78.600 63.200 ;
        RECT 47.800 62.800 78.600 63.100 ;
        RECT 101.400 63.100 101.800 63.200 ;
        RECT 103.800 63.100 104.200 63.200 ;
        RECT 101.400 62.800 104.200 63.100 ;
        RECT 137.400 63.100 137.800 63.200 ;
        RECT 154.200 63.100 154.600 63.200 ;
        RECT 137.400 62.800 154.600 63.100 ;
        RECT 63.800 62.100 64.200 62.200 ;
        RECT 71.800 62.100 72.200 62.200 ;
        RECT 89.400 62.100 89.800 62.200 ;
        RECT 63.800 61.800 89.800 62.100 ;
        RECT 121.400 62.100 121.800 62.200 ;
        RECT 142.200 62.100 142.600 62.200 ;
        RECT 121.400 61.800 142.600 62.100 ;
        RECT 143.000 62.100 143.400 62.200 ;
        RECT 144.600 62.100 145.000 62.200 ;
        RECT 143.000 61.800 145.000 62.100 ;
        RECT 170.200 62.100 170.600 62.200 ;
        RECT 171.000 62.100 171.400 62.200 ;
        RECT 170.200 61.800 171.400 62.100 ;
        RECT 79.800 61.100 80.200 61.200 ;
        RECT 83.800 61.100 84.200 61.200 ;
        RECT 79.800 60.800 84.200 61.100 ;
        RECT 85.400 61.100 85.800 61.200 ;
        RECT 131.000 61.100 131.400 61.200 ;
        RECT 85.400 60.800 131.400 61.100 ;
        RECT 165.400 61.100 165.800 61.200 ;
        RECT 169.400 61.100 169.800 61.200 ;
        RECT 165.400 60.800 169.800 61.100 ;
        RECT 47.000 60.100 47.400 60.200 ;
        RECT 52.600 60.100 53.000 60.200 ;
        RECT 47.000 59.800 53.000 60.100 ;
        RECT 77.400 60.100 77.800 60.200 ;
        RECT 83.800 60.100 84.200 60.200 ;
        RECT 98.200 60.100 98.600 60.200 ;
        RECT 77.400 59.800 98.600 60.100 ;
        RECT 100.600 60.100 101.000 60.200 ;
        RECT 101.400 60.100 101.800 60.200 ;
        RECT 110.200 60.100 110.600 60.200 ;
        RECT 100.600 59.800 110.600 60.100 ;
        RECT 123.800 60.100 124.200 60.200 ;
        RECT 136.600 60.100 137.000 60.200 ;
        RECT 123.800 59.800 137.000 60.100 ;
        RECT 142.200 60.100 142.600 60.200 ;
        RECT 151.800 60.100 152.200 60.200 ;
        RECT 142.200 59.800 152.200 60.100 ;
        RECT 161.400 60.100 161.800 60.200 ;
        RECT 163.800 60.100 164.200 60.200 ;
        RECT 161.400 59.800 164.200 60.100 ;
        RECT 9.400 59.100 9.800 59.200 ;
        RECT 20.600 59.100 21.000 59.200 ;
        RECT 23.800 59.100 24.200 59.200 ;
        RECT 67.000 59.100 67.400 59.200 ;
        RECT 118.200 59.100 118.600 59.200 ;
        RECT 157.400 59.100 157.800 59.200 ;
        RECT 166.200 59.100 166.600 59.200 ;
        RECT 9.400 58.800 118.600 59.100 ;
        RECT 119.000 58.800 166.600 59.100 ;
        RECT 171.000 59.100 171.400 59.200 ;
        RECT 176.600 59.100 177.000 59.200 ;
        RECT 171.000 58.800 177.000 59.100 ;
        RECT 119.000 58.200 119.300 58.800 ;
        RECT 44.600 57.800 45.000 58.200 ;
        RECT 100.600 57.800 101.000 58.200 ;
        RECT 119.000 57.800 119.400 58.200 ;
        RECT 132.600 58.100 133.000 58.200 ;
        RECT 142.200 58.100 142.600 58.200 ;
        RECT 132.600 57.800 142.600 58.100 ;
        RECT 147.800 58.100 148.200 58.200 ;
        RECT 159.800 58.100 160.200 58.200 ;
        RECT 147.800 57.800 160.200 58.100 ;
        RECT 179.000 57.800 179.400 58.200 ;
        RECT 4.600 57.100 5.000 57.200 ;
        RECT 22.200 57.100 22.600 57.200 ;
        RECT 4.600 56.800 22.600 57.100 ;
        RECT 27.800 56.800 28.200 57.200 ;
        RECT 44.600 57.100 44.900 57.800 ;
        RECT 100.600 57.200 100.900 57.800 ;
        RECT 179.000 57.200 179.300 57.800 ;
        RECT 46.200 57.100 46.600 57.200 ;
        RECT 44.600 56.800 46.600 57.100 ;
        RECT 100.600 56.800 101.000 57.200 ;
        RECT 115.000 57.100 115.400 57.200 ;
        RECT 149.400 57.100 149.800 57.200 ;
        RECT 157.400 57.100 157.800 57.200 ;
        RECT 168.600 57.100 169.000 57.200 ;
        RECT 115.000 56.800 169.000 57.100 ;
        RECT 179.000 56.800 179.400 57.200 ;
        RECT 7.000 56.100 7.400 56.200 ;
        RECT 13.400 56.100 13.800 56.200 ;
        RECT 24.600 56.100 25.000 56.200 ;
        RECT 7.000 55.800 25.000 56.100 ;
        RECT 27.800 56.100 28.100 56.800 ;
        RECT 33.400 56.100 33.800 56.200 ;
        RECT 27.800 55.800 33.800 56.100 ;
        RECT 49.400 56.100 49.800 56.200 ;
        RECT 50.200 56.100 50.600 56.200 ;
        RECT 49.400 55.800 50.600 56.100 ;
        RECT 55.800 56.100 56.200 56.200 ;
        RECT 58.200 56.100 58.600 56.200 ;
        RECT 62.200 56.100 62.600 56.200 ;
        RECT 55.800 55.800 62.600 56.100 ;
        RECT 73.400 56.100 73.800 56.200 ;
        RECT 91.800 56.100 92.200 56.200 ;
        RECT 73.400 55.800 92.200 56.100 ;
        RECT 119.000 55.800 119.400 56.200 ;
        RECT 133.400 56.100 133.800 56.200 ;
        RECT 139.000 56.100 139.400 56.200 ;
        RECT 143.000 56.100 143.400 56.200 ;
        RECT 133.400 55.800 136.100 56.100 ;
        RECT 139.000 55.800 143.400 56.100 ;
        RECT 143.800 56.100 144.200 56.200 ;
        RECT 163.800 56.100 164.200 56.200 ;
        RECT 165.400 56.100 165.800 56.200 ;
        RECT 143.800 55.800 165.800 56.100 ;
        RECT 170.200 56.100 170.600 56.200 ;
        RECT 179.800 56.100 180.200 56.200 ;
        RECT 170.200 55.800 180.200 56.100 ;
        RECT 119.000 55.200 119.300 55.800 ;
        RECT 2.200 55.100 2.600 55.200 ;
        RECT 5.400 55.100 5.800 55.200 ;
        RECT 2.200 54.800 5.800 55.100 ;
        RECT 22.200 54.800 22.600 55.200 ;
        RECT 26.200 55.100 26.600 55.200 ;
        RECT 28.600 55.100 29.000 55.200 ;
        RECT 26.200 54.800 29.000 55.100 ;
        RECT 30.200 55.100 30.600 55.200 ;
        RECT 40.600 55.100 41.000 55.200 ;
        RECT 30.200 54.800 41.000 55.100 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 49.400 55.100 49.800 55.200 ;
        RECT 47.000 54.800 49.800 55.100 ;
        RECT 51.800 55.100 52.200 55.200 ;
        RECT 54.200 55.100 54.600 55.200 ;
        RECT 56.600 55.100 57.000 55.200 ;
        RECT 51.800 54.800 57.000 55.100 ;
        RECT 70.200 54.800 70.600 55.200 ;
        RECT 78.200 55.100 78.600 55.200 ;
        RECT 94.200 55.100 94.600 55.200 ;
        RECT 78.200 54.800 94.600 55.100 ;
        RECT 97.400 55.100 97.800 55.200 ;
        RECT 99.000 55.100 99.400 55.200 ;
        RECT 111.800 55.100 112.200 55.200 ;
        RECT 97.400 54.800 99.400 55.100 ;
        RECT 106.200 54.800 112.200 55.100 ;
        RECT 113.400 55.100 113.800 55.200 ;
        RECT 114.200 55.100 114.600 55.200 ;
        RECT 113.400 54.800 114.600 55.100 ;
        RECT 119.000 54.800 119.400 55.200 ;
        RECT 120.600 55.100 121.000 55.200 ;
        RECT 130.200 55.100 130.600 55.200 ;
        RECT 120.600 54.800 130.600 55.100 ;
        RECT 135.000 54.800 135.400 55.200 ;
        RECT 135.800 55.100 136.100 55.800 ;
        RECT 138.200 55.100 138.600 55.200 ;
        RECT 135.800 54.800 138.600 55.100 ;
        RECT 140.600 55.100 141.000 55.200 ;
        RECT 141.400 55.100 141.800 55.200 ;
        RECT 140.600 54.800 141.800 55.100 ;
        RECT 155.800 55.100 156.200 55.200 ;
        RECT 158.200 55.100 158.600 55.200 ;
        RECT 155.800 54.800 158.600 55.100 ;
        RECT 176.600 54.800 177.000 55.200 ;
        RECT 22.200 54.200 22.500 54.800 ;
        RECT 70.200 54.200 70.500 54.800 ;
        RECT 106.200 54.700 106.600 54.800 ;
        RECT 3.000 53.800 3.400 54.200 ;
        RECT 22.200 53.800 22.600 54.200 ;
        RECT 24.600 54.100 25.000 54.200 ;
        RECT 40.600 54.100 41.000 54.200 ;
        RECT 67.800 54.100 68.200 54.200 ;
        RECT 24.600 53.800 68.200 54.100 ;
        RECT 70.200 53.800 70.600 54.200 ;
        RECT 81.400 54.100 81.800 54.200 ;
        RECT 82.200 54.100 82.600 54.200 ;
        RECT 81.400 53.800 82.600 54.100 ;
        RECT 96.600 54.100 97.000 54.200 ;
        RECT 99.800 54.100 100.200 54.200 ;
        RECT 96.600 53.800 100.200 54.100 ;
        RECT 123.800 54.100 124.200 54.200 ;
        RECT 124.600 54.100 125.000 54.200 ;
        RECT 123.800 53.800 125.000 54.100 ;
        RECT 135.000 54.100 135.300 54.800 ;
        RECT 176.600 54.200 176.900 54.800 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 149.400 54.100 149.800 54.200 ;
        RECT 155.800 54.100 156.200 54.200 ;
        RECT 135.000 53.800 145.700 54.100 ;
        RECT 149.400 53.800 156.200 54.100 ;
        RECT 161.400 54.100 161.800 54.200 ;
        RECT 168.600 54.100 169.000 54.200 ;
        RECT 161.400 53.800 169.000 54.100 ;
        RECT 176.600 53.800 177.000 54.200 ;
        RECT 3.000 53.200 3.300 53.800 ;
        RECT 145.400 53.200 145.700 53.800 ;
        RECT 3.000 52.800 3.400 53.200 ;
        RECT 6.200 53.100 6.600 53.200 ;
        RECT 16.600 53.100 17.000 53.200 ;
        RECT 21.400 53.100 21.800 53.200 ;
        RECT 31.800 53.100 32.200 53.200 ;
        RECT 6.200 52.800 32.200 53.100 ;
        RECT 48.600 53.100 49.000 53.200 ;
        RECT 50.200 53.100 50.600 53.200 ;
        RECT 48.600 52.800 50.600 53.100 ;
        RECT 51.000 53.100 51.400 53.200 ;
        RECT 61.400 53.100 61.800 53.200 ;
        RECT 51.000 52.800 61.800 53.100 ;
        RECT 67.000 53.100 67.400 53.200 ;
        RECT 69.400 53.100 69.800 53.200 ;
        RECT 67.000 52.800 69.800 53.100 ;
        RECT 73.400 53.100 73.800 53.200 ;
        RECT 75.800 53.100 76.200 53.200 ;
        RECT 73.400 52.800 76.200 53.100 ;
        RECT 90.200 53.100 90.600 53.200 ;
        RECT 97.400 53.100 97.800 53.200 ;
        RECT 90.200 52.800 97.800 53.100 ;
        RECT 145.400 52.800 145.800 53.200 ;
        RECT 55.800 52.100 56.200 52.200 ;
        RECT 62.200 52.100 62.600 52.200 ;
        RECT 55.800 51.800 62.600 52.100 ;
        RECT 64.600 52.100 65.000 52.200 ;
        RECT 79.000 52.100 79.400 52.200 ;
        RECT 80.600 52.100 81.000 52.200 ;
        RECT 87.000 52.100 87.400 52.200 ;
        RECT 64.600 51.800 87.400 52.100 ;
        RECT 87.800 52.100 88.200 52.200 ;
        RECT 105.400 52.100 105.800 52.200 ;
        RECT 110.200 52.100 110.600 52.200 ;
        RECT 87.800 51.800 110.600 52.100 ;
        RECT 127.800 52.100 128.200 52.200 ;
        RECT 136.600 52.100 137.000 52.200 ;
        RECT 127.800 51.800 137.000 52.100 ;
        RECT 154.200 52.100 154.600 52.200 ;
        RECT 175.000 52.100 175.400 52.200 ;
        RECT 154.200 51.800 175.400 52.100 ;
        RECT 17.400 51.100 17.800 51.200 ;
        RECT 19.800 51.100 20.200 51.200 ;
        RECT 44.600 51.100 45.000 51.200 ;
        RECT 17.400 50.800 45.000 51.100 ;
        RECT 103.000 51.100 103.400 51.200 ;
        RECT 116.600 51.100 117.000 51.200 ;
        RECT 103.000 50.800 117.000 51.100 ;
        RECT 119.800 51.100 120.200 51.200 ;
        RECT 143.800 51.100 144.200 51.200 ;
        RECT 119.800 50.800 144.200 51.100 ;
        RECT 153.400 51.100 153.800 51.200 ;
        RECT 155.000 51.100 155.400 51.200 ;
        RECT 153.400 50.800 155.400 51.100 ;
        RECT 156.600 51.100 157.000 51.200 ;
        RECT 161.400 51.100 161.800 51.200 ;
        RECT 156.600 50.800 161.800 51.100 ;
        RECT 173.400 51.100 173.800 51.200 ;
        RECT 177.400 51.100 177.800 51.200 ;
        RECT 173.400 50.800 177.800 51.100 ;
        RECT 9.400 49.800 9.800 50.200 ;
        RECT 41.400 50.100 41.800 50.200 ;
        RECT 45.400 50.100 45.800 50.200 ;
        RECT 53.400 50.100 53.800 50.200 ;
        RECT 41.400 49.800 53.800 50.100 ;
        RECT 91.800 50.100 92.200 50.200 ;
        RECT 107.800 50.100 108.200 50.200 ;
        RECT 91.800 49.800 108.200 50.100 ;
        RECT 118.200 50.100 118.600 50.200 ;
        RECT 122.200 50.100 122.600 50.200 ;
        RECT 118.200 49.800 122.600 50.100 ;
        RECT 156.600 49.800 157.000 50.200 ;
        RECT 7.800 49.100 8.200 49.200 ;
        RECT 9.400 49.100 9.700 49.800 ;
        RECT 7.800 48.800 9.700 49.100 ;
        RECT 35.000 49.100 35.400 49.200 ;
        RECT 43.800 49.100 44.200 49.200 ;
        RECT 44.600 49.100 45.000 49.200 ;
        RECT 35.000 48.800 45.000 49.100 ;
        RECT 59.800 49.100 60.200 49.200 ;
        RECT 67.800 49.100 68.200 49.200 ;
        RECT 68.600 49.100 69.000 49.200 ;
        RECT 59.800 48.800 69.000 49.100 ;
        RECT 91.000 49.100 91.400 49.200 ;
        RECT 97.400 49.100 97.800 49.200 ;
        RECT 109.400 49.100 109.800 49.200 ;
        RECT 121.400 49.100 121.800 49.200 ;
        RECT 123.800 49.100 124.200 49.200 ;
        RECT 91.000 48.800 97.800 49.100 ;
        RECT 108.600 48.800 124.200 49.100 ;
        RECT 155.800 49.100 156.200 49.200 ;
        RECT 156.600 49.100 156.900 49.800 ;
        RECT 155.800 48.800 156.900 49.100 ;
        RECT 166.200 49.100 166.600 49.200 ;
        RECT 167.800 49.100 168.200 49.200 ;
        RECT 166.200 48.800 168.200 49.100 ;
        RECT 16.600 47.800 17.000 48.200 ;
        RECT 61.400 48.100 61.800 48.200 ;
        RECT 71.800 48.100 72.200 48.200 ;
        RECT 61.400 47.800 72.200 48.100 ;
        RECT 75.000 48.100 75.400 48.200 ;
        RECT 92.600 48.100 93.000 48.200 ;
        RECT 75.000 47.800 93.000 48.100 ;
        RECT 98.200 48.100 98.600 48.200 ;
        RECT 101.400 48.100 101.800 48.200 ;
        RECT 98.200 47.800 101.800 48.100 ;
        RECT 104.600 48.100 105.000 48.200 ;
        RECT 108.600 48.100 109.000 48.200 ;
        RECT 119.800 48.100 120.200 48.200 ;
        RECT 104.600 47.800 120.200 48.100 ;
        RECT 120.600 48.100 121.000 48.200 ;
        RECT 136.600 48.100 137.000 48.200 ;
        RECT 120.600 47.800 137.000 48.100 ;
        RECT 146.200 48.100 146.600 48.200 ;
        RECT 159.800 48.100 160.200 48.200 ;
        RECT 146.200 47.800 160.200 48.100 ;
        RECT 166.200 47.800 166.600 48.200 ;
        RECT 168.600 47.800 169.000 48.200 ;
        RECT 12.600 47.100 13.000 47.200 ;
        RECT 16.600 47.100 16.900 47.800 ;
        RECT 166.200 47.200 166.500 47.800 ;
        RECT 168.600 47.200 168.900 47.800 ;
        RECT 12.600 46.800 16.900 47.100 ;
        RECT 27.800 46.800 28.200 47.200 ;
        RECT 38.200 46.800 38.600 47.200 ;
        RECT 52.600 47.100 53.000 47.200 ;
        RECT 54.200 47.100 54.600 47.200 ;
        RECT 55.000 47.100 55.400 47.200 ;
        RECT 52.600 46.800 53.700 47.100 ;
        RECT 54.200 46.800 55.400 47.100 ;
        RECT 65.400 47.100 65.800 47.200 ;
        RECT 68.600 47.100 69.000 47.200 ;
        RECT 65.400 46.800 69.000 47.100 ;
        RECT 76.600 47.100 77.000 47.200 ;
        RECT 83.800 47.100 84.200 47.200 ;
        RECT 93.400 47.100 93.800 47.200 ;
        RECT 76.600 46.800 81.700 47.100 ;
        RECT 83.800 46.800 93.800 47.100 ;
        RECT 112.600 47.100 113.000 47.200 ;
        RECT 127.800 47.100 128.200 47.200 ;
        RECT 112.600 46.800 128.200 47.100 ;
        RECT 131.000 47.100 131.400 47.200 ;
        RECT 133.400 47.100 133.800 47.200 ;
        RECT 131.000 46.800 133.800 47.100 ;
        RECT 134.200 46.800 134.600 47.200 ;
        RECT 159.800 46.800 160.200 47.200 ;
        RECT 166.200 46.800 166.600 47.200 ;
        RECT 168.600 46.800 169.000 47.200 ;
        RECT 27.800 46.200 28.100 46.800 ;
        RECT 16.600 46.100 17.000 46.200 ;
        RECT 23.000 46.100 23.400 46.200 ;
        RECT 27.800 46.100 28.200 46.200 ;
        RECT 16.600 45.800 28.200 46.100 ;
        RECT 31.800 46.100 32.200 46.200 ;
        RECT 38.200 46.100 38.500 46.800 ;
        RECT 31.800 45.800 38.500 46.100 ;
        RECT 53.400 46.100 53.700 46.800 ;
        RECT 81.400 46.200 81.700 46.800 ;
        RECT 59.800 46.100 60.200 46.200 ;
        RECT 63.000 46.100 63.400 46.200 ;
        RECT 53.400 45.800 63.400 46.100 ;
        RECT 81.400 45.800 81.800 46.200 ;
        RECT 87.000 46.100 87.400 46.200 ;
        RECT 97.400 46.100 97.800 46.200 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 87.000 45.800 103.400 46.100 ;
        RECT 112.600 46.100 113.000 46.200 ;
        RECT 122.200 46.100 122.600 46.200 ;
        RECT 112.600 45.800 122.600 46.100 ;
        RECT 123.800 46.100 124.200 46.200 ;
        RECT 127.000 46.100 127.400 46.200 ;
        RECT 123.800 45.800 127.400 46.100 ;
        RECT 128.600 46.100 129.000 46.200 ;
        RECT 134.200 46.100 134.500 46.800 ;
        RECT 128.600 45.800 134.500 46.100 ;
        RECT 150.200 46.100 150.600 46.200 ;
        RECT 159.800 46.100 160.100 46.800 ;
        RECT 169.400 46.100 169.800 46.200 ;
        RECT 150.200 45.800 169.800 46.100 ;
        RECT 171.800 46.100 172.200 46.200 ;
        RECT 175.800 46.100 176.200 46.200 ;
        RECT 171.800 45.800 176.200 46.100 ;
        RECT 8.600 45.100 9.000 45.200 ;
        RECT 19.000 45.100 19.400 45.200 ;
        RECT 8.600 44.800 19.400 45.100 ;
        RECT 42.200 45.100 42.600 45.200 ;
        RECT 71.800 45.100 72.200 45.200 ;
        RECT 42.200 44.800 72.200 45.100 ;
        RECT 81.400 45.100 81.800 45.200 ;
        RECT 82.200 45.100 82.600 45.200 ;
        RECT 81.400 44.800 82.600 45.100 ;
        RECT 116.600 45.100 117.000 45.200 ;
        RECT 118.200 45.100 118.600 45.200 ;
        RECT 116.600 44.800 118.600 45.100 ;
        RECT 120.600 45.100 121.000 45.200 ;
        RECT 124.600 45.100 125.000 45.200 ;
        RECT 120.600 44.800 125.000 45.100 ;
        RECT 154.200 45.100 154.600 45.200 ;
        RECT 155.000 45.100 155.400 45.200 ;
        RECT 167.000 45.100 167.400 45.200 ;
        RECT 154.200 44.800 167.400 45.100 ;
        RECT 169.400 45.100 169.800 45.200 ;
        RECT 174.200 45.100 174.600 45.200 ;
        RECT 169.400 44.800 174.600 45.100 ;
        RECT 176.600 44.800 177.000 45.200 ;
        RECT 176.600 44.200 176.900 44.800 ;
        RECT 15.000 44.100 15.400 44.200 ;
        RECT 25.400 44.100 25.800 44.200 ;
        RECT 35.800 44.100 36.200 44.200 ;
        RECT 57.400 44.100 57.800 44.200 ;
        RECT 15.000 43.800 57.800 44.100 ;
        RECT 87.800 44.100 88.200 44.200 ;
        RECT 89.400 44.100 89.800 44.200 ;
        RECT 87.800 43.800 89.800 44.100 ;
        RECT 136.600 44.100 137.000 44.200 ;
        RECT 146.200 44.100 146.600 44.200 ;
        RECT 136.600 43.800 146.600 44.100 ;
        RECT 155.800 44.100 156.200 44.200 ;
        RECT 158.200 44.100 158.600 44.200 ;
        RECT 155.800 43.800 158.600 44.100 ;
        RECT 176.600 43.800 177.000 44.200 ;
        RECT 20.600 43.100 21.000 43.200 ;
        RECT 81.400 43.100 81.800 43.200 ;
        RECT 100.600 43.100 101.000 43.200 ;
        RECT 104.600 43.100 105.000 43.200 ;
        RECT 114.200 43.100 114.600 43.200 ;
        RECT 20.600 42.800 80.900 43.100 ;
        RECT 81.400 42.800 114.600 43.100 ;
        RECT 19.800 42.100 20.200 42.200 ;
        RECT 28.600 42.100 29.000 42.200 ;
        RECT 78.200 42.100 78.600 42.200 ;
        RECT 19.800 41.800 78.600 42.100 ;
        RECT 80.600 42.100 80.900 42.800 ;
        RECT 148.600 42.100 149.000 42.200 ;
        RECT 162.200 42.100 162.600 42.200 ;
        RECT 80.600 41.800 162.600 42.100 ;
        RECT 171.800 41.800 172.200 42.200 ;
        RECT 171.800 41.200 172.100 41.800 ;
        RECT 160.600 41.100 161.000 41.200 ;
        RECT 163.000 41.100 163.400 41.200 ;
        RECT 164.600 41.100 165.000 41.200 ;
        RECT 160.600 40.800 165.000 41.100 ;
        RECT 171.800 40.800 172.200 41.200 ;
        RECT 14.200 40.100 14.600 40.200 ;
        RECT 20.600 40.100 21.000 40.200 ;
        RECT 14.200 39.800 21.000 40.100 ;
        RECT 44.600 40.100 45.000 40.200 ;
        RECT 53.400 40.100 53.800 40.200 ;
        RECT 44.600 39.800 53.800 40.100 ;
        RECT 97.400 40.100 97.800 40.200 ;
        RECT 101.400 40.100 101.800 40.200 ;
        RECT 97.400 39.800 101.800 40.100 ;
        RECT 151.800 40.100 152.200 40.200 ;
        RECT 158.200 40.100 158.600 40.200 ;
        RECT 167.000 40.100 167.400 40.200 ;
        RECT 151.800 39.800 167.400 40.100 ;
        RECT 171.800 40.100 172.200 40.200 ;
        RECT 172.600 40.100 173.000 40.200 ;
        RECT 171.800 39.800 173.000 40.100 ;
        RECT 70.200 39.100 70.600 39.200 ;
        RECT 80.600 39.100 81.000 39.200 ;
        RECT 65.400 38.800 81.000 39.100 ;
        RECT 94.200 39.100 94.600 39.200 ;
        RECT 99.000 39.100 99.400 39.200 ;
        RECT 103.000 39.100 103.400 39.200 ;
        RECT 94.200 38.800 103.400 39.100 ;
        RECT 140.600 39.100 141.000 39.200 ;
        RECT 141.400 39.100 141.800 39.200 ;
        RECT 140.600 38.800 141.800 39.100 ;
        RECT 65.400 38.200 65.700 38.800 ;
        RECT 65.400 37.800 65.800 38.200 ;
        RECT 79.000 38.100 79.400 38.200 ;
        RECT 106.200 38.100 106.600 38.200 ;
        RECT 79.000 37.800 106.600 38.100 ;
        RECT 28.600 37.100 29.000 37.200 ;
        RECT 34.200 37.100 34.600 37.200 ;
        RECT 46.200 37.100 46.600 37.200 ;
        RECT 28.600 36.800 46.600 37.100 ;
        RECT 48.600 37.100 49.000 37.200 ;
        RECT 51.000 37.100 51.400 37.200 ;
        RECT 48.600 36.800 51.400 37.100 ;
        RECT 54.200 36.800 54.600 37.200 ;
        RECT 55.000 37.100 55.400 37.200 ;
        RECT 55.800 37.100 56.200 37.200 ;
        RECT 55.000 36.800 56.200 37.100 ;
        RECT 76.600 37.100 77.000 37.200 ;
        RECT 88.600 37.100 89.000 37.200 ;
        RECT 91.800 37.100 92.200 37.200 ;
        RECT 76.600 36.800 84.100 37.100 ;
        RECT 88.600 36.800 92.200 37.100 ;
        RECT 104.600 37.100 105.000 37.200 ;
        RECT 109.400 37.100 109.800 37.200 ;
        RECT 104.600 36.800 109.800 37.100 ;
        RECT 174.200 37.100 174.600 37.200 ;
        RECT 178.200 37.100 178.600 37.200 ;
        RECT 174.200 36.800 178.600 37.100 ;
        RECT 3.800 36.100 4.200 36.200 ;
        RECT 13.400 36.100 13.800 36.200 ;
        RECT 3.800 35.800 13.800 36.100 ;
        RECT 18.200 35.800 18.600 36.200 ;
        RECT 27.800 36.100 28.200 36.200 ;
        RECT 28.600 36.100 29.000 36.200 ;
        RECT 35.000 36.100 35.400 36.200 ;
        RECT 27.800 35.800 35.400 36.100 ;
        RECT 40.600 36.100 41.000 36.200 ;
        RECT 54.200 36.100 54.500 36.800 ;
        RECT 83.800 36.200 84.100 36.800 ;
        RECT 40.600 35.800 54.500 36.100 ;
        RECT 55.000 36.100 55.400 36.200 ;
        RECT 55.800 36.100 56.200 36.200 ;
        RECT 55.000 35.800 56.200 36.100 ;
        RECT 64.600 36.100 65.000 36.200 ;
        RECT 65.400 36.100 65.800 36.200 ;
        RECT 67.800 36.100 68.200 36.200 ;
        RECT 64.600 35.800 68.200 36.100 ;
        RECT 82.200 36.100 82.600 36.200 ;
        RECT 83.000 36.100 83.400 36.200 ;
        RECT 82.200 35.800 83.400 36.100 ;
        RECT 83.800 35.800 84.200 36.200 ;
        RECT 97.400 36.100 97.800 36.200 ;
        RECT 91.000 35.800 97.800 36.100 ;
        RECT 100.600 36.100 101.000 36.200 ;
        RECT 163.800 36.100 164.200 36.200 ;
        RECT 100.600 35.800 164.200 36.100 ;
        RECT 175.800 35.800 176.200 36.200 ;
        RECT 4.600 35.100 5.000 35.200 ;
        RECT 10.200 35.100 10.600 35.200 ;
        RECT 4.600 34.800 10.600 35.100 ;
        RECT 18.200 35.100 18.500 35.800 ;
        RECT 91.000 35.200 91.300 35.800 ;
        RECT 23.000 35.100 23.400 35.200 ;
        RECT 58.200 35.100 58.600 35.200 ;
        RECT 71.800 35.100 72.200 35.200 ;
        RECT 18.200 34.800 58.600 35.100 ;
        RECT 69.400 34.800 72.200 35.100 ;
        RECT 77.400 35.100 77.800 35.200 ;
        RECT 82.200 35.100 82.600 35.200 ;
        RECT 84.600 35.100 85.000 35.200 ;
        RECT 77.400 34.800 85.000 35.100 ;
        RECT 91.000 34.800 91.400 35.200 ;
        RECT 95.800 34.800 96.200 35.200 ;
        RECT 107.000 35.100 107.400 35.200 ;
        RECT 115.800 35.100 116.200 35.200 ;
        RECT 119.800 35.100 120.200 35.200 ;
        RECT 107.000 34.800 115.300 35.100 ;
        RECT 115.800 34.800 120.200 35.100 ;
        RECT 122.200 35.100 122.600 35.200 ;
        RECT 123.000 35.100 123.400 35.200 ;
        RECT 122.200 34.800 123.400 35.100 ;
        RECT 161.400 35.100 161.800 35.200 ;
        RECT 170.200 35.100 170.600 35.200 ;
        RECT 161.400 34.800 170.600 35.100 ;
        RECT 175.000 35.100 175.400 35.200 ;
        RECT 175.800 35.100 176.100 35.800 ;
        RECT 175.000 34.800 176.100 35.100 ;
        RECT 69.400 34.200 69.700 34.800 ;
        RECT 22.200 34.100 22.600 34.200 ;
        RECT 30.200 34.100 30.600 34.200 ;
        RECT 22.200 33.800 30.600 34.100 ;
        RECT 42.200 33.800 42.600 34.200 ;
        RECT 47.000 34.100 47.400 34.200 ;
        RECT 50.200 34.100 50.600 34.200 ;
        RECT 47.000 33.800 52.900 34.100 ;
        RECT 69.400 33.800 69.800 34.200 ;
        RECT 87.800 34.100 88.200 34.200 ;
        RECT 95.800 34.100 96.100 34.800 ;
        RECT 87.800 33.800 96.100 34.100 ;
        RECT 106.200 34.100 106.600 34.200 ;
        RECT 108.600 34.100 109.000 34.200 ;
        RECT 106.200 33.800 109.000 34.100 ;
        RECT 115.000 34.100 115.300 34.800 ;
        RECT 118.200 34.100 118.600 34.200 ;
        RECT 120.600 34.100 121.000 34.200 ;
        RECT 115.000 33.800 121.000 34.100 ;
        RECT 127.000 34.100 127.400 34.200 ;
        RECT 167.800 34.100 168.200 34.200 ;
        RECT 170.200 34.100 170.600 34.200 ;
        RECT 127.000 33.800 134.500 34.100 ;
        RECT 167.800 33.800 170.600 34.100 ;
        RECT 171.000 33.800 171.400 34.200 ;
        RECT 3.000 33.100 3.400 33.200 ;
        RECT 29.400 33.100 29.800 33.200 ;
        RECT 31.800 33.100 32.200 33.200 ;
        RECT 35.000 33.100 35.400 33.200 ;
        RECT 3.000 32.800 35.400 33.100 ;
        RECT 36.600 33.100 37.000 33.200 ;
        RECT 42.200 33.100 42.500 33.800 ;
        RECT 52.600 33.200 52.900 33.800 ;
        RECT 134.200 33.200 134.500 33.800 ;
        RECT 171.000 33.200 171.300 33.800 ;
        RECT 49.400 33.100 49.800 33.200 ;
        RECT 36.600 32.800 49.800 33.100 ;
        RECT 52.600 32.800 53.000 33.200 ;
        RECT 53.400 33.100 53.800 33.200 ;
        RECT 59.800 33.100 60.200 33.200 ;
        RECT 68.600 33.100 69.000 33.200 ;
        RECT 75.800 33.100 76.200 33.200 ;
        RECT 53.400 32.800 76.200 33.100 ;
        RECT 79.800 33.100 80.200 33.200 ;
        RECT 81.400 33.100 81.800 33.200 ;
        RECT 79.800 32.800 81.800 33.100 ;
        RECT 87.000 33.100 87.400 33.200 ;
        RECT 103.800 33.100 104.200 33.200 ;
        RECT 114.200 33.100 114.600 33.200 ;
        RECT 87.000 32.800 104.200 33.100 ;
        RECT 107.800 32.800 114.600 33.100 ;
        RECT 122.200 33.100 122.600 33.200 ;
        RECT 123.000 33.100 123.400 33.200 ;
        RECT 122.200 32.800 123.400 33.100 ;
        RECT 134.200 32.800 134.600 33.200 ;
        RECT 171.000 32.800 171.400 33.200 ;
        RECT 107.800 32.200 108.100 32.800 ;
        RECT 19.000 32.100 19.400 32.200 ;
        RECT 43.800 32.100 44.200 32.200 ;
        RECT 19.000 31.800 44.200 32.100 ;
        RECT 53.400 32.100 53.800 32.200 ;
        RECT 63.000 32.100 63.400 32.200 ;
        RECT 53.400 31.800 63.400 32.100 ;
        RECT 63.800 32.100 64.200 32.200 ;
        RECT 69.400 32.100 69.800 32.200 ;
        RECT 63.800 31.800 69.800 32.100 ;
        RECT 75.800 32.100 76.200 32.200 ;
        RECT 85.400 32.100 85.800 32.200 ;
        RECT 99.000 32.100 99.400 32.200 ;
        RECT 75.800 31.800 99.400 32.100 ;
        RECT 107.800 31.800 108.200 32.200 ;
        RECT 123.000 32.100 123.400 32.200 ;
        RECT 137.400 32.100 137.800 32.200 ;
        RECT 139.000 32.100 139.400 32.200 ;
        RECT 147.000 32.100 147.400 32.200 ;
        RECT 153.400 32.100 153.800 32.200 ;
        RECT 123.000 31.800 153.800 32.100 ;
        RECT 159.000 32.100 159.400 32.200 ;
        RECT 164.600 32.100 165.000 32.200 ;
        RECT 159.000 31.800 165.000 32.100 ;
        RECT 107.800 31.100 108.200 31.200 ;
        RECT 116.600 31.100 117.000 31.200 ;
        RECT 123.800 31.100 124.200 31.200 ;
        RECT 107.800 30.800 124.200 31.100 ;
        RECT 125.400 31.100 125.800 31.200 ;
        RECT 143.000 31.100 143.400 31.200 ;
        RECT 125.400 30.800 143.400 31.100 ;
        RECT 9.400 30.100 9.800 30.200 ;
        RECT 17.400 30.100 17.800 30.200 ;
        RECT 9.400 29.800 17.800 30.100 ;
        RECT 65.400 30.100 65.800 30.200 ;
        RECT 74.200 30.100 74.600 30.200 ;
        RECT 65.400 29.800 74.600 30.100 ;
        RECT 169.400 30.100 169.800 30.200 ;
        RECT 171.000 30.100 171.400 30.200 ;
        RECT 169.400 29.800 171.400 30.100 ;
        RECT 6.200 29.100 6.600 29.200 ;
        RECT 18.200 29.100 18.600 29.200 ;
        RECT 21.400 29.100 21.800 29.200 ;
        RECT 28.600 29.100 29.000 29.200 ;
        RECT 6.200 28.800 29.000 29.100 ;
        RECT 31.000 29.100 31.400 29.200 ;
        RECT 37.400 29.100 37.800 29.200 ;
        RECT 31.000 28.800 37.800 29.100 ;
        RECT 55.000 29.100 55.400 29.200 ;
        RECT 64.600 29.100 65.000 29.200 ;
        RECT 55.000 28.800 65.000 29.100 ;
        RECT 67.800 29.100 68.200 29.200 ;
        RECT 79.800 29.100 80.200 29.200 ;
        RECT 67.800 28.800 80.200 29.100 ;
        RECT 82.200 29.100 82.600 29.200 ;
        RECT 83.000 29.100 83.400 29.200 ;
        RECT 91.800 29.100 92.200 29.200 ;
        RECT 82.200 28.800 92.200 29.100 ;
        RECT 92.600 29.100 93.000 29.200 ;
        RECT 100.600 29.100 101.000 29.200 ;
        RECT 92.600 28.800 101.000 29.100 ;
        RECT 119.000 29.100 119.400 29.200 ;
        RECT 130.200 29.100 130.600 29.200 ;
        RECT 119.000 28.800 130.600 29.100 ;
        RECT 143.800 29.100 144.200 29.200 ;
        RECT 144.600 29.100 145.000 29.200 ;
        RECT 179.800 29.100 180.200 29.200 ;
        RECT 143.800 28.800 145.000 29.100 ;
        RECT 169.400 28.800 180.200 29.100 ;
        RECT 169.400 28.200 169.700 28.800 ;
        RECT 15.800 28.100 16.200 28.200 ;
        RECT 17.400 28.100 17.800 28.200 ;
        RECT 43.000 28.100 43.400 28.200 ;
        RECT 15.800 27.800 43.400 28.100 ;
        RECT 124.600 28.100 125.000 28.200 ;
        RECT 126.200 28.100 126.600 28.200 ;
        RECT 124.600 27.800 126.600 28.100 ;
        RECT 169.400 28.100 169.800 28.200 ;
        RECT 170.200 28.100 170.600 28.200 ;
        RECT 169.400 27.800 170.600 28.100 ;
        RECT 12.600 27.100 13.000 27.200 ;
        RECT 15.000 27.100 15.400 27.200 ;
        RECT 12.600 26.800 15.400 27.100 ;
        RECT 15.800 27.100 16.200 27.200 ;
        RECT 27.800 27.100 28.200 27.200 ;
        RECT 15.800 26.800 28.200 27.100 ;
        RECT 43.000 27.100 43.400 27.200 ;
        RECT 45.400 27.100 45.800 27.200 ;
        RECT 61.400 27.100 61.800 27.200 ;
        RECT 43.000 26.800 61.800 27.100 ;
        RECT 76.600 27.100 77.000 27.200 ;
        RECT 79.800 27.100 80.200 27.200 ;
        RECT 76.600 26.800 80.200 27.100 ;
        RECT 88.600 27.100 89.000 27.200 ;
        RECT 95.800 27.100 96.200 27.200 ;
        RECT 88.600 26.800 96.200 27.100 ;
        RECT 121.400 27.100 121.800 27.200 ;
        RECT 132.600 27.100 133.000 27.200 ;
        RECT 121.400 26.800 133.000 27.100 ;
        RECT 153.400 27.100 153.800 27.200 ;
        RECT 173.400 27.100 173.800 27.200 ;
        RECT 153.400 26.800 173.800 27.100 ;
        RECT 4.600 26.100 5.000 26.200 ;
        RECT 11.800 26.100 12.200 26.200 ;
        RECT 4.600 25.800 12.200 26.100 ;
        RECT 20.600 26.100 21.000 26.200 ;
        RECT 40.600 26.100 41.000 26.200 ;
        RECT 20.600 25.800 41.000 26.100 ;
        RECT 48.600 26.100 49.000 26.200 ;
        RECT 51.000 26.100 51.400 26.200 ;
        RECT 55.000 26.100 55.400 26.200 ;
        RECT 48.600 25.800 55.400 26.100 ;
        RECT 63.800 26.100 64.200 26.200 ;
        RECT 74.200 26.100 74.600 26.200 ;
        RECT 97.400 26.100 97.800 26.200 ;
        RECT 98.200 26.100 98.600 26.200 ;
        RECT 63.800 25.800 98.600 26.100 ;
        RECT 103.800 26.100 104.200 26.200 ;
        RECT 111.000 26.100 111.400 26.200 ;
        RECT 103.800 25.800 111.400 26.100 ;
        RECT 114.200 26.100 114.600 26.200 ;
        RECT 115.800 26.100 116.200 26.200 ;
        RECT 127.000 26.100 127.400 26.200 ;
        RECT 150.200 26.100 150.600 26.200 ;
        RECT 158.200 26.100 158.600 26.200 ;
        RECT 161.400 26.100 161.800 26.200 ;
        RECT 114.200 25.800 161.800 26.100 ;
        RECT 174.200 26.100 174.600 26.200 ;
        RECT 179.000 26.100 179.400 26.200 ;
        RECT 174.200 25.800 179.400 26.100 ;
        RECT 130.200 25.200 130.500 25.800 ;
        RECT 3.000 25.100 3.400 25.200 ;
        RECT 3.800 25.100 4.200 25.200 ;
        RECT 3.000 24.800 4.200 25.100 ;
        RECT 13.400 25.100 13.800 25.200 ;
        RECT 15.000 25.100 15.400 25.200 ;
        RECT 23.000 25.100 23.400 25.200 ;
        RECT 13.400 24.800 23.400 25.100 ;
        RECT 42.200 24.800 42.600 25.200 ;
        RECT 46.200 25.100 46.600 25.200 ;
        RECT 49.400 25.100 49.800 25.200 ;
        RECT 67.800 25.100 68.200 25.200 ;
        RECT 46.200 24.800 68.200 25.100 ;
        RECT 114.200 25.100 114.600 25.200 ;
        RECT 116.600 25.100 117.000 25.200 ;
        RECT 123.800 25.100 124.200 25.200 ;
        RECT 114.200 24.800 124.200 25.100 ;
        RECT 130.200 24.800 130.600 25.200 ;
        RECT 136.600 24.800 137.000 25.200 ;
        RECT 146.200 25.100 146.600 25.200 ;
        RECT 151.000 25.100 151.400 25.200 ;
        RECT 146.200 24.800 151.400 25.100 ;
        RECT 154.200 25.100 154.600 25.200 ;
        RECT 173.400 25.100 173.800 25.200 ;
        RECT 154.200 24.800 173.800 25.100 ;
        RECT 42.200 24.100 42.500 24.800 ;
        RECT 136.600 24.200 136.900 24.800 ;
        RECT 60.600 24.100 61.000 24.200 ;
        RECT 75.000 24.100 75.400 24.200 ;
        RECT 42.200 23.800 49.700 24.100 ;
        RECT 60.600 23.800 75.400 24.100 ;
        RECT 136.600 23.800 137.000 24.200 ;
        RECT 168.600 24.100 169.000 24.200 ;
        RECT 171.800 24.100 172.200 24.200 ;
        RECT 168.600 23.800 172.200 24.100 ;
        RECT 49.400 23.200 49.700 23.800 ;
        RECT 49.400 22.800 49.800 23.200 ;
        RECT 50.200 23.100 50.600 23.200 ;
        RECT 61.400 23.100 61.800 23.200 ;
        RECT 50.200 22.800 61.800 23.100 ;
        RECT 84.600 23.100 85.000 23.200 ;
        RECT 137.400 23.100 137.800 23.200 ;
        RECT 141.400 23.100 141.800 23.200 ;
        RECT 156.600 23.100 157.000 23.200 ;
        RECT 169.400 23.100 169.800 23.200 ;
        RECT 84.600 22.800 169.800 23.100 ;
        RECT 171.800 23.100 172.200 23.200 ;
        RECT 174.200 23.100 174.600 23.200 ;
        RECT 171.800 22.800 174.600 23.100 ;
        RECT 34.200 22.100 34.600 22.200 ;
        RECT 37.400 22.100 37.800 22.200 ;
        RECT 50.200 22.100 50.600 22.200 ;
        RECT 51.000 22.100 51.400 22.200 ;
        RECT 34.200 21.800 37.800 22.100 ;
        RECT 49.400 21.800 51.400 22.100 ;
        RECT 51.800 22.100 52.200 22.200 ;
        RECT 68.600 22.100 69.000 22.200 ;
        RECT 51.800 21.800 69.000 22.100 ;
        RECT 136.600 22.100 137.000 22.200 ;
        RECT 145.400 22.100 145.800 22.200 ;
        RECT 136.600 21.800 145.800 22.100 ;
        RECT 169.400 22.100 169.800 22.200 ;
        RECT 178.200 22.100 178.600 22.200 ;
        RECT 169.400 21.800 178.600 22.100 ;
        RECT 96.600 21.100 97.000 21.200 ;
        RECT 99.800 21.100 100.200 21.200 ;
        RECT 112.600 21.100 113.000 21.200 ;
        RECT 118.200 21.100 118.600 21.200 ;
        RECT 121.400 21.100 121.800 21.200 ;
        RECT 96.600 20.800 121.800 21.100 ;
        RECT 75.000 20.100 75.400 20.200 ;
        RECT 87.800 20.100 88.200 20.200 ;
        RECT 111.800 20.100 112.200 20.200 ;
        RECT 75.000 19.800 112.200 20.100 ;
        RECT 162.200 19.800 162.600 20.200 ;
        RECT 37.400 19.100 37.800 19.200 ;
        RECT 41.400 19.100 41.800 19.200 ;
        RECT 37.400 18.800 41.800 19.100 ;
        RECT 79.800 19.100 80.200 19.200 ;
        RECT 80.600 19.100 81.000 19.200 ;
        RECT 91.000 19.100 91.400 19.200 ;
        RECT 79.800 18.800 91.400 19.100 ;
        RECT 97.400 19.100 97.800 19.200 ;
        RECT 98.200 19.100 98.600 19.200 ;
        RECT 107.000 19.100 107.400 19.200 ;
        RECT 97.400 18.800 107.400 19.100 ;
        RECT 159.800 19.100 160.200 19.200 ;
        RECT 162.200 19.100 162.500 19.800 ;
        RECT 159.800 18.800 162.500 19.100 ;
        RECT 9.400 18.100 9.800 18.200 ;
        RECT 19.000 18.100 19.400 18.200 ;
        RECT 9.400 17.800 19.400 18.100 ;
        RECT 136.600 17.800 137.000 18.200 ;
        RECT 140.600 18.100 141.000 18.200 ;
        RECT 152.600 18.100 153.000 18.200 ;
        RECT 159.000 18.100 159.400 18.200 ;
        RECT 140.600 17.800 159.400 18.100 ;
        RECT 136.600 17.200 136.900 17.800 ;
        RECT 4.600 17.100 5.000 17.200 ;
        RECT 22.200 17.100 22.600 17.200 ;
        RECT 4.600 16.800 22.600 17.100 ;
        RECT 27.800 17.100 28.200 17.200 ;
        RECT 67.000 17.100 67.400 17.200 ;
        RECT 27.800 16.800 67.400 17.100 ;
        RECT 87.800 17.100 88.200 17.200 ;
        RECT 100.600 17.100 101.000 17.200 ;
        RECT 87.800 16.800 101.000 17.100 ;
        RECT 110.200 16.800 110.600 17.200 ;
        RECT 136.600 16.800 137.000 17.200 ;
        RECT 140.600 17.100 141.000 17.200 ;
        RECT 147.000 17.100 147.400 17.200 ;
        RECT 148.600 17.100 149.000 17.200 ;
        RECT 179.000 17.100 179.400 17.200 ;
        RECT 140.600 16.800 149.000 17.100 ;
        RECT 155.000 16.800 179.400 17.100 ;
        RECT 1.400 16.100 1.800 16.200 ;
        RECT 5.400 16.100 5.800 16.200 ;
        RECT 1.400 15.800 5.800 16.100 ;
        RECT 31.800 16.100 32.200 16.200 ;
        RECT 60.600 16.100 61.000 16.200 ;
        RECT 31.800 15.800 61.000 16.100 ;
        RECT 68.600 16.100 69.000 16.200 ;
        RECT 79.000 16.100 79.400 16.200 ;
        RECT 68.600 15.800 79.400 16.100 ;
        RECT 86.200 15.800 86.600 16.200 ;
        RECT 95.000 16.100 95.400 16.200 ;
        RECT 95.800 16.100 96.200 16.200 ;
        RECT 95.000 15.800 96.200 16.100 ;
        RECT 103.800 16.100 104.200 16.200 ;
        RECT 110.200 16.100 110.500 16.800 ;
        RECT 103.800 15.800 110.500 16.100 ;
        RECT 114.200 16.100 114.600 16.200 ;
        RECT 115.800 16.100 116.200 16.200 ;
        RECT 114.200 15.800 116.200 16.100 ;
        RECT 117.400 16.100 117.800 16.200 ;
        RECT 119.800 16.100 120.200 16.200 ;
        RECT 117.400 15.800 120.200 16.100 ;
        RECT 122.200 16.100 122.600 16.200 ;
        RECT 128.600 16.100 129.000 16.200 ;
        RECT 122.200 15.800 129.000 16.100 ;
        RECT 148.600 16.100 149.000 16.200 ;
        RECT 155.000 16.100 155.300 16.800 ;
        RECT 148.600 15.800 155.300 16.100 ;
        RECT 155.800 15.800 156.200 16.200 ;
        RECT 166.200 16.100 166.600 16.200 ;
        RECT 170.200 16.100 170.600 16.200 ;
        RECT 166.200 15.800 170.600 16.100 ;
        RECT 172.600 16.100 173.000 16.200 ;
        RECT 175.800 16.100 176.200 16.200 ;
        RECT 172.600 15.800 176.200 16.100 ;
        RECT 3.800 15.100 4.200 15.200 ;
        RECT 6.200 15.100 6.600 15.200 ;
        RECT 3.800 14.800 6.600 15.100 ;
        RECT 7.800 15.100 8.200 15.200 ;
        RECT 11.000 15.100 11.400 15.200 ;
        RECT 20.600 15.100 21.000 15.200 ;
        RECT 7.800 14.800 21.000 15.100 ;
        RECT 22.200 15.100 22.600 15.200 ;
        RECT 39.000 15.100 39.400 15.200 ;
        RECT 22.200 14.800 39.400 15.100 ;
        RECT 41.400 15.100 41.800 15.200 ;
        RECT 51.000 15.100 51.400 15.200 ;
        RECT 65.400 15.100 65.800 15.200 ;
        RECT 75.000 15.100 75.400 15.200 ;
        RECT 41.400 14.800 75.400 15.100 ;
        RECT 86.200 15.100 86.500 15.800 ;
        RECT 92.600 15.100 93.000 15.200 ;
        RECT 86.200 14.800 93.000 15.100 ;
        RECT 95.000 15.100 95.400 15.200 ;
        RECT 109.400 15.100 109.800 15.200 ;
        RECT 117.400 15.100 117.800 15.200 ;
        RECT 95.000 14.800 117.800 15.100 ;
        RECT 120.600 15.100 121.000 15.200 ;
        RECT 123.800 15.100 124.200 15.200 ;
        RECT 120.600 14.800 124.200 15.100 ;
        RECT 130.200 15.100 130.600 15.200 ;
        RECT 138.200 15.100 138.600 15.200 ;
        RECT 130.200 14.800 138.600 15.100 ;
        RECT 143.000 15.100 143.400 15.200 ;
        RECT 148.600 15.100 148.900 15.800 ;
        RECT 143.000 14.800 148.900 15.100 ;
        RECT 151.800 15.100 152.200 15.200 ;
        RECT 155.800 15.100 156.100 15.800 ;
        RECT 151.800 14.800 156.100 15.100 ;
        RECT 164.600 15.100 165.000 15.200 ;
        RECT 177.400 15.100 177.800 15.200 ;
        RECT 178.200 15.100 178.600 15.200 ;
        RECT 164.600 14.800 178.600 15.100 ;
        RECT 31.800 14.100 32.200 14.200 ;
        RECT 41.400 14.100 41.800 14.200 ;
        RECT 31.800 13.800 41.800 14.100 ;
        RECT 49.400 13.800 49.800 14.200 ;
        RECT 52.600 14.100 53.000 14.200 ;
        RECT 53.400 14.100 53.800 14.200 ;
        RECT 52.600 13.800 53.800 14.100 ;
        RECT 55.800 13.800 56.200 14.200 ;
        RECT 57.400 14.100 57.800 14.200 ;
        RECT 59.000 14.100 59.400 14.200 ;
        RECT 71.800 14.100 72.200 14.200 ;
        RECT 73.400 14.100 73.800 14.200 ;
        RECT 115.000 14.100 115.400 14.200 ;
        RECT 57.400 13.800 115.400 14.100 ;
        RECT 146.200 14.100 146.600 14.200 ;
        RECT 147.800 14.100 148.200 14.200 ;
        RECT 163.000 14.100 163.400 14.200 ;
        RECT 146.200 13.800 163.400 14.100 ;
        RECT 170.200 13.800 170.600 14.200 ;
        RECT 12.600 13.100 13.000 13.200 ;
        RECT 16.600 13.100 17.000 13.200 ;
        RECT 12.600 12.800 17.000 13.100 ;
        RECT 37.400 13.100 37.800 13.200 ;
        RECT 44.600 13.100 45.000 13.200 ;
        RECT 37.400 12.800 45.000 13.100 ;
        RECT 49.400 13.100 49.700 13.800 ;
        RECT 55.800 13.100 56.100 13.800 ;
        RECT 170.200 13.200 170.500 13.800 ;
        RECT 49.400 12.800 56.100 13.100 ;
        RECT 56.600 13.100 57.000 13.200 ;
        RECT 59.800 13.100 60.200 13.200 ;
        RECT 56.600 12.800 60.200 13.100 ;
        RECT 117.400 13.100 117.800 13.200 ;
        RECT 119.000 13.100 119.400 13.200 ;
        RECT 119.800 13.100 120.200 13.200 ;
        RECT 117.400 12.800 120.200 13.100 ;
        RECT 140.600 13.100 141.000 13.200 ;
        RECT 144.600 13.100 145.000 13.200 ;
        RECT 149.400 13.100 149.800 13.200 ;
        RECT 140.600 12.800 149.800 13.100 ;
        RECT 170.200 12.800 170.600 13.200 ;
        RECT 19.000 12.100 19.400 12.200 ;
        RECT 21.400 12.100 21.800 12.200 ;
        RECT 19.000 11.800 21.800 12.100 ;
        RECT 112.600 12.100 113.000 12.200 ;
        RECT 123.800 12.100 124.200 12.200 ;
        RECT 112.600 11.800 124.200 12.100 ;
        RECT 19.800 11.100 20.200 11.200 ;
        RECT 23.000 11.100 23.400 11.200 ;
        RECT 19.800 10.800 23.400 11.100 ;
        RECT 122.200 11.100 122.600 11.200 ;
        RECT 123.000 11.100 123.400 11.200 ;
        RECT 122.200 10.800 123.400 11.100 ;
        RECT 163.800 11.100 164.200 11.200 ;
        RECT 176.600 11.100 177.000 11.200 ;
        RECT 163.800 10.800 177.000 11.100 ;
        RECT 9.400 9.800 9.800 10.200 ;
        RECT 16.600 10.100 17.000 10.200 ;
        RECT 19.000 10.100 19.400 10.200 ;
        RECT 16.600 9.800 19.400 10.100 ;
        RECT 96.600 10.100 97.000 10.200 ;
        RECT 113.400 10.100 113.800 10.200 ;
        RECT 96.600 9.800 113.800 10.100 ;
        RECT 169.400 10.100 169.800 10.200 ;
        RECT 171.800 10.100 172.200 10.200 ;
        RECT 169.400 9.800 172.200 10.100 ;
        RECT 179.000 9.800 179.400 10.200 ;
        RECT 6.200 9.100 6.600 9.200 ;
        RECT 9.400 9.100 9.700 9.800 ;
        RECT 179.000 9.200 179.300 9.800 ;
        RECT 6.200 8.800 9.700 9.100 ;
        RECT 27.800 9.100 28.200 9.200 ;
        RECT 33.400 9.100 33.800 9.200 ;
        RECT 27.800 8.800 33.800 9.100 ;
        RECT 49.400 8.800 49.800 9.200 ;
        RECT 66.200 9.100 66.600 9.200 ;
        RECT 69.400 9.100 69.800 9.200 ;
        RECT 66.200 8.800 69.800 9.100 ;
        RECT 104.600 9.100 105.000 9.200 ;
        RECT 111.800 9.100 112.200 9.200 ;
        RECT 127.000 9.100 127.400 9.200 ;
        RECT 104.600 8.800 127.400 9.100 ;
        RECT 138.200 8.800 138.600 9.200 ;
        RECT 151.000 9.100 151.400 9.200 ;
        RECT 160.600 9.100 161.000 9.200 ;
        RECT 167.800 9.100 168.200 9.200 ;
        RECT 151.000 8.800 168.200 9.100 ;
        RECT 179.000 8.800 179.400 9.200 ;
        RECT 11.000 7.800 11.400 8.200 ;
        RECT 15.800 8.100 16.200 8.200 ;
        RECT 22.200 8.100 22.600 8.200 ;
        RECT 15.800 7.800 22.600 8.100 ;
        RECT 37.400 7.800 37.800 8.200 ;
        RECT 41.400 8.100 41.800 8.200 ;
        RECT 49.400 8.100 49.700 8.800 ;
        RECT 41.400 7.800 49.700 8.100 ;
        RECT 52.600 7.800 53.000 8.200 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 129.400 8.100 129.800 8.200 ;
        RECT 130.200 8.100 130.600 8.200 ;
        RECT 129.400 7.800 130.600 8.100 ;
        RECT 135.800 8.100 136.200 8.200 ;
        RECT 138.200 8.100 138.500 8.800 ;
        RECT 135.800 7.800 138.500 8.100 ;
        RECT 139.800 8.100 140.200 8.200 ;
        RECT 140.600 8.100 141.000 8.200 ;
        RECT 139.800 7.800 141.000 8.100 ;
        RECT 171.000 7.800 171.400 8.200 ;
        RECT 5.400 7.100 5.800 7.200 ;
        RECT 11.000 7.100 11.300 7.800 ;
        RECT 5.400 6.800 11.300 7.100 ;
        RECT 12.600 6.800 13.000 7.200 ;
        RECT 24.600 7.100 25.000 7.200 ;
        RECT 27.800 7.100 28.200 7.200 ;
        RECT 24.600 6.800 28.200 7.100 ;
        RECT 29.400 7.100 29.800 7.200 ;
        RECT 37.400 7.100 37.700 7.800 ;
        RECT 52.600 7.100 52.900 7.800 ;
        RECT 29.400 6.800 52.900 7.100 ;
        RECT 71.800 6.800 72.200 7.200 ;
        RECT 78.200 7.100 78.500 7.800 ;
        RECT 171.000 7.200 171.300 7.800 ;
        RECT 83.000 7.100 83.400 7.200 ;
        RECT 78.200 6.800 83.400 7.100 ;
        RECT 90.200 7.100 90.600 7.200 ;
        RECT 146.200 7.100 146.600 7.200 ;
        RECT 90.200 6.800 146.600 7.100 ;
        RECT 149.400 7.100 149.800 7.200 ;
        RECT 153.400 7.100 153.800 7.200 ;
        RECT 149.400 6.800 153.800 7.100 ;
        RECT 171.000 6.800 171.400 7.200 ;
        RECT 172.600 6.800 173.000 7.200 ;
        RECT 8.600 6.100 9.000 6.200 ;
        RECT 12.600 6.100 12.900 6.800 ;
        RECT 8.600 5.800 12.900 6.100 ;
        RECT 20.600 6.100 21.000 6.200 ;
        RECT 23.800 6.100 24.200 6.200 ;
        RECT 26.200 6.100 26.600 6.200 ;
        RECT 47.000 6.100 47.400 6.200 ;
        RECT 50.200 6.100 50.600 6.200 ;
        RECT 20.600 5.800 50.600 6.100 ;
        RECT 55.800 6.100 56.200 6.200 ;
        RECT 63.000 6.100 63.400 6.200 ;
        RECT 55.800 5.800 63.400 6.100 ;
        RECT 71.800 6.100 72.100 6.800 ;
        RECT 73.400 6.100 73.800 6.200 ;
        RECT 71.800 5.800 73.800 6.100 ;
        RECT 77.400 6.100 77.800 6.200 ;
        RECT 86.200 6.100 86.600 6.200 ;
        RECT 93.400 6.100 93.800 6.200 ;
        RECT 77.400 5.800 86.600 6.100 ;
        RECT 89.400 5.800 93.800 6.100 ;
        RECT 102.200 6.100 102.600 6.300 ;
        RECT 172.600 6.200 172.900 6.800 ;
        RECT 116.600 6.100 117.000 6.200 ;
        RECT 102.200 5.800 117.000 6.100 ;
        RECT 122.200 6.100 122.600 6.200 ;
        RECT 143.800 6.100 144.200 6.200 ;
        RECT 122.200 5.800 144.200 6.100 ;
        RECT 150.200 6.100 150.600 6.200 ;
        RECT 151.000 6.100 151.400 6.200 ;
        RECT 150.200 5.800 151.400 6.100 ;
        RECT 172.600 5.800 173.000 6.200 ;
        RECT 89.400 5.200 89.700 5.800 ;
        RECT 19.800 5.100 20.200 5.200 ;
        RECT 89.400 5.100 89.800 5.200 ;
        RECT 19.800 4.800 89.800 5.100 ;
        RECT 98.200 5.100 98.600 5.200 ;
        RECT 147.000 5.100 147.400 5.200 ;
        RECT 98.200 4.800 147.400 5.100 ;
      LAYER via3 ;
        RECT 51.800 168.800 52.200 169.200 ;
        RECT 40.600 165.800 41.000 166.200 ;
        RECT 103.800 165.800 104.200 166.200 ;
        RECT 93.400 164.800 93.800 165.200 ;
        RECT 44.600 163.800 45.000 164.200 ;
        RECT 101.400 163.800 101.800 164.200 ;
        RECT 174.200 163.800 174.600 164.200 ;
        RECT 169.400 161.800 169.800 162.200 ;
        RECT 87.800 157.800 88.200 158.200 ;
        RECT 59.800 155.800 60.200 156.200 ;
        RECT 173.400 155.800 173.800 156.200 ;
        RECT 172.600 151.800 173.000 152.200 ;
        RECT 87.000 149.800 87.400 150.200 ;
        RECT 158.200 147.800 158.600 148.200 ;
        RECT 93.400 146.800 93.800 147.200 ;
        RECT 103.000 146.800 103.400 147.200 ;
        RECT 155.800 146.800 156.200 147.200 ;
        RECT 157.400 146.800 157.800 147.200 ;
        RECT 77.400 145.800 77.800 146.200 ;
        RECT 100.600 145.800 101.000 146.200 ;
        RECT 45.400 144.800 45.800 145.200 ;
        RECT 69.400 140.800 69.800 141.200 ;
        RECT 59.800 138.800 60.200 139.200 ;
        RECT 64.600 136.800 65.000 137.200 ;
        RECT 103.800 136.800 104.200 137.200 ;
        RECT 23.000 135.800 23.400 136.200 ;
        RECT 31.000 135.800 31.400 136.200 ;
        RECT 59.800 135.800 60.200 136.200 ;
        RECT 34.200 134.800 34.600 135.200 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 53.400 133.800 53.800 134.200 ;
        RECT 56.600 133.800 57.000 134.200 ;
        RECT 103.000 133.800 103.400 134.200 ;
        RECT 41.400 132.800 41.800 133.200 ;
        RECT 83.000 132.800 83.400 133.200 ;
        RECT 132.600 132.800 133.000 133.200 ;
        RECT 168.600 132.800 169.000 133.200 ;
        RECT 6.200 131.800 6.600 132.200 ;
        RECT 166.200 130.800 166.600 131.200 ;
        RECT 28.600 124.800 29.000 125.200 ;
        RECT 63.800 124.800 64.200 125.200 ;
        RECT 161.400 124.800 161.800 125.200 ;
        RECT 15.800 123.800 16.200 124.200 ;
        RECT 39.800 123.800 40.200 124.200 ;
        RECT 64.600 123.800 65.000 124.200 ;
        RECT 115.000 122.800 115.400 123.200 ;
        RECT 97.400 120.800 97.800 121.200 ;
        RECT 171.800 117.800 172.200 118.200 ;
        RECT 47.800 115.800 48.200 116.200 ;
        RECT 157.400 115.800 157.800 116.200 ;
        RECT 72.600 114.800 73.000 115.200 ;
        RECT 85.400 114.800 85.800 115.200 ;
        RECT 160.600 114.800 161.000 115.200 ;
        RECT 107.000 113.800 107.400 114.200 ;
        RECT 31.000 111.800 31.400 112.200 ;
        RECT 151.800 111.800 152.200 112.200 ;
        RECT 42.200 106.800 42.600 107.200 ;
        RECT 78.200 106.800 78.600 107.200 ;
        RECT 83.800 106.800 84.200 107.200 ;
        RECT 147.000 106.800 147.400 107.200 ;
        RECT 167.800 105.800 168.200 106.200 ;
        RECT 41.400 103.800 41.800 104.200 ;
        RECT 113.400 101.800 113.800 102.200 ;
        RECT 129.400 101.800 129.800 102.200 ;
        RECT 76.600 100.800 77.000 101.200 ;
        RECT 98.200 100.800 98.600 101.200 ;
        RECT 163.000 100.800 163.400 101.200 ;
        RECT 42.200 98.800 42.600 99.200 ;
        RECT 164.600 98.800 165.000 99.200 ;
        RECT 39.800 96.800 40.200 97.200 ;
        RECT 47.000 95.800 47.400 96.200 ;
        RECT 59.800 94.800 60.200 95.200 ;
        RECT 113.400 94.800 113.800 95.200 ;
        RECT 159.000 94.800 159.400 95.200 ;
        RECT 19.800 93.800 20.200 94.200 ;
        RECT 55.800 92.800 56.200 93.200 ;
        RECT 42.200 91.800 42.600 92.200 ;
        RECT 46.200 91.800 46.600 92.200 ;
        RECT 129.400 90.800 129.800 91.200 ;
        RECT 102.200 89.800 102.600 90.200 ;
        RECT 115.000 88.800 115.400 89.200 ;
        RECT 163.800 88.800 164.200 89.200 ;
        RECT 67.800 87.800 68.200 88.200 ;
        RECT 93.400 87.800 93.800 88.200 ;
        RECT 173.400 87.800 173.800 88.200 ;
        RECT 22.200 86.800 22.600 87.200 ;
        RECT 159.800 86.800 160.200 87.200 ;
        RECT 23.800 85.800 24.200 86.200 ;
        RECT 34.200 85.800 34.600 86.200 ;
        RECT 43.800 85.800 44.200 86.200 ;
        RECT 98.200 85.800 98.600 86.200 ;
        RECT 171.000 85.800 171.400 86.200 ;
        RECT 19.000 84.800 19.400 85.200 ;
        RECT 155.000 84.800 155.400 85.200 ;
        RECT 45.400 83.800 45.800 84.200 ;
        RECT 175.000 83.800 175.400 84.200 ;
        RECT 75.000 82.800 75.400 83.200 ;
        RECT 132.600 79.800 133.000 80.200 ;
        RECT 28.600 77.800 29.000 78.200 ;
        RECT 86.200 77.800 86.600 78.200 ;
        RECT 63.800 76.800 64.200 77.200 ;
        RECT 87.000 76.800 87.400 77.200 ;
        RECT 111.800 76.800 112.200 77.200 ;
        RECT 23.000 75.800 23.400 76.200 ;
        RECT 49.400 75.800 49.800 76.200 ;
        RECT 114.200 74.800 114.600 75.200 ;
        RECT 128.600 74.800 129.000 75.200 ;
        RECT 133.400 74.800 133.800 75.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 143.800 73.800 144.200 74.200 ;
        RECT 174.200 73.800 174.600 74.200 ;
        RECT 116.600 72.800 117.000 73.200 ;
        RECT 140.600 72.800 141.000 73.200 ;
        RECT 117.400 71.800 117.800 72.200 ;
        RECT 175.800 71.800 176.200 72.200 ;
        RECT 153.400 70.800 153.800 71.200 ;
        RECT 86.200 68.800 86.600 69.200 ;
        RECT 156.600 68.800 157.000 69.200 ;
        RECT 56.600 67.800 57.000 68.200 ;
        RECT 161.400 67.800 161.800 68.200 ;
        RECT 91.800 66.800 92.200 67.200 ;
        RECT 99.800 66.800 100.200 67.200 ;
        RECT 20.600 64.800 21.000 65.200 ;
        RECT 83.000 64.800 83.400 65.200 ;
        RECT 168.600 64.800 169.000 65.200 ;
        RECT 72.600 63.800 73.000 64.200 ;
        RECT 95.800 63.800 96.200 64.200 ;
        RECT 78.200 62.800 78.600 63.200 ;
        RECT 142.200 61.800 142.600 62.200 ;
        RECT 171.000 61.800 171.400 62.200 ;
        RECT 101.400 59.800 101.800 60.200 ;
        RECT 166.200 58.800 166.600 59.200 ;
        RECT 176.600 58.800 177.000 59.200 ;
        RECT 163.800 55.800 164.200 56.200 ;
        RECT 179.800 55.800 180.200 56.200 ;
        RECT 158.200 54.800 158.600 55.200 ;
        RECT 40.600 53.800 41.000 54.200 ;
        RECT 82.200 53.800 82.600 54.200 ;
        RECT 124.600 53.800 125.000 54.200 ;
        RECT 87.000 51.800 87.400 52.200 ;
        RECT 44.600 48.800 45.000 49.200 ;
        RECT 67.800 48.800 68.200 49.200 ;
        RECT 167.800 48.800 168.200 49.200 ;
        RECT 119.800 47.800 120.200 48.200 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 82.200 44.800 82.600 45.200 ;
        RECT 124.600 44.800 125.000 45.200 ;
        RECT 155.000 44.800 155.400 45.200 ;
        RECT 167.000 44.800 167.400 45.200 ;
        RECT 146.200 43.800 146.600 44.200 ;
        RECT 114.200 42.800 114.600 43.200 ;
        RECT 53.400 39.800 53.800 40.200 ;
        RECT 172.600 39.800 173.000 40.200 ;
        RECT 70.200 38.800 70.600 39.200 ;
        RECT 55.800 36.800 56.200 37.200 ;
        RECT 178.200 36.800 178.600 37.200 ;
        RECT 55.800 35.800 56.200 36.200 ;
        RECT 23.000 34.800 23.400 35.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 123.000 34.800 123.400 35.200 ;
        RECT 118.200 33.800 118.600 34.200 ;
        RECT 31.800 32.800 32.200 33.200 ;
        RECT 35.000 32.800 35.400 33.200 ;
        RECT 123.000 32.800 123.400 33.200 ;
        RECT 63.000 31.800 63.400 32.200 ;
        RECT 99.000 31.800 99.400 32.200 ;
        RECT 116.600 30.800 117.000 31.200 ;
        RECT 74.200 29.800 74.600 30.200 ;
        RECT 171.000 29.800 171.400 30.200 ;
        RECT 170.200 27.800 170.600 28.200 ;
        RECT 27.800 26.800 28.200 27.200 ;
        RECT 98.200 25.800 98.600 26.200 ;
        RECT 49.400 24.800 49.800 25.200 ;
        RECT 169.400 22.800 169.800 23.200 ;
        RECT 87.800 19.800 88.200 20.200 ;
        RECT 115.800 15.800 116.200 16.200 ;
        RECT 119.800 15.800 120.200 16.200 ;
        RECT 128.600 15.800 129.000 16.200 ;
        RECT 178.200 14.800 178.600 15.200 ;
        RECT 53.400 13.800 53.800 14.200 ;
        RECT 119.800 12.800 120.200 13.200 ;
        RECT 130.200 7.800 130.600 8.200 ;
        RECT 151.000 5.800 151.400 6.200 ;
      LAYER metal4 ;
        RECT 51.800 168.800 52.200 169.200 ;
        RECT 6.200 165.800 6.600 166.200 ;
        RECT 40.600 165.800 41.000 166.200 ;
        RECT 6.200 132.200 6.500 165.800 ;
        RECT 40.600 155.200 40.900 165.800 ;
        RECT 44.600 163.800 45.000 164.200 ;
        RECT 40.600 154.800 41.000 155.200 ;
        RECT 15.000 154.100 15.400 154.200 ;
        RECT 15.000 153.800 16.100 154.100 ;
        RECT 6.200 131.800 6.600 132.200 ;
        RECT 15.800 124.200 16.100 153.800 ;
        RECT 23.000 136.100 23.400 136.200 ;
        RECT 22.200 135.800 23.400 136.100 ;
        RECT 31.000 135.800 31.400 136.200 ;
        RECT 15.800 123.800 16.200 124.200 ;
        RECT 22.200 106.200 22.500 135.800 ;
        RECT 28.600 124.800 29.000 125.200 ;
        RECT 25.400 116.800 25.800 117.200 ;
        RECT 22.200 105.800 22.600 106.200 ;
        RECT 19.000 97.800 19.400 98.200 ;
        RECT 19.000 85.200 19.300 97.800 ;
        RECT 19.800 93.800 20.200 94.200 ;
        RECT 19.000 84.800 19.400 85.200 ;
        RECT 19.800 65.100 20.100 93.800 ;
        RECT 22.200 86.800 22.600 87.200 ;
        RECT 20.600 65.100 21.000 65.200 ;
        RECT 19.800 64.800 21.000 65.100 ;
        RECT 3.000 52.800 3.400 53.200 ;
        RECT 3.000 33.200 3.300 52.800 ;
        RECT 19.800 42.200 20.100 64.800 ;
        RECT 22.200 54.200 22.500 86.800 ;
        RECT 25.400 86.200 25.700 116.800 ;
        RECT 23.800 86.100 24.200 86.200 ;
        RECT 24.600 86.100 25.000 86.200 ;
        RECT 23.800 85.800 25.000 86.100 ;
        RECT 25.400 85.800 25.800 86.200 ;
        RECT 27.800 81.800 28.200 82.200 ;
        RECT 23.000 75.800 23.400 76.200 ;
        RECT 22.200 53.800 22.600 54.200 ;
        RECT 19.800 41.800 20.200 42.200 ;
        RECT 23.000 35.200 23.300 75.800 ;
        RECT 27.800 46.200 28.100 81.800 ;
        RECT 28.600 78.200 28.900 124.800 ;
        RECT 31.000 112.200 31.300 135.800 ;
        RECT 34.200 135.100 34.600 135.200 ;
        RECT 33.400 134.800 34.600 135.100 ;
        RECT 31.000 111.800 31.400 112.200 ;
        RECT 33.400 96.200 33.700 134.800 ;
        RECT 34.200 134.200 34.500 134.800 ;
        RECT 34.200 133.800 34.600 134.200 ;
        RECT 41.400 133.100 41.800 133.200 ;
        RECT 42.200 133.100 42.600 133.200 ;
        RECT 41.400 132.800 42.600 133.100 ;
        RECT 44.600 132.200 44.900 163.800 ;
        RECT 45.400 146.800 45.800 147.200 ;
        RECT 48.600 147.100 49.000 147.200 ;
        RECT 49.400 147.100 49.800 147.200 ;
        RECT 48.600 146.800 49.800 147.100 ;
        RECT 45.400 145.200 45.700 146.800 ;
        RECT 45.400 144.800 45.800 145.200 ;
        RECT 46.200 144.800 46.600 145.200 ;
        RECT 44.600 131.800 45.000 132.200 ;
        RECT 45.400 129.800 45.800 130.200 ;
        RECT 39.800 123.800 40.200 124.200 ;
        RECT 35.000 112.800 35.400 113.200 ;
        RECT 33.400 95.800 33.800 96.200 ;
        RECT 33.400 86.100 33.800 86.200 ;
        RECT 34.200 86.100 34.600 86.200 ;
        RECT 33.400 85.800 34.600 86.100 ;
        RECT 28.600 77.800 29.000 78.200 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 27.800 36.100 28.200 36.200 ;
        RECT 28.600 36.100 28.900 77.800 ;
        RECT 27.800 35.800 28.900 36.100 ;
        RECT 23.000 34.800 23.400 35.200 ;
        RECT 3.000 32.800 3.400 33.200 ;
        RECT 3.000 25.200 3.300 32.800 ;
        RECT 27.800 27.200 28.100 35.800 ;
        RECT 35.000 33.200 35.300 112.800 ;
        RECT 39.800 97.200 40.100 123.800 ;
        RECT 43.000 107.800 43.400 108.200 ;
        RECT 42.200 106.800 42.600 107.200 ;
        RECT 41.400 104.100 41.800 104.200 ;
        RECT 40.600 103.800 41.800 104.100 ;
        RECT 39.800 96.800 40.200 97.200 ;
        RECT 40.600 54.200 40.900 103.800 ;
        RECT 42.200 101.200 42.500 106.800 ;
        RECT 42.200 100.800 42.600 101.200 ;
        RECT 42.200 99.200 42.500 100.800 ;
        RECT 42.200 98.800 42.600 99.200 ;
        RECT 42.200 91.800 42.600 92.200 ;
        RECT 40.600 53.800 41.000 54.200 ;
        RECT 42.200 45.200 42.500 91.800 ;
        RECT 43.000 87.200 43.300 107.800 ;
        RECT 45.400 98.200 45.700 129.800 ;
        RECT 46.200 103.200 46.500 144.800 ;
        RECT 51.800 142.200 52.100 168.800 ;
        RECT 103.800 165.800 104.200 166.200 ;
        RECT 159.000 165.800 159.400 166.200 ;
        RECT 164.600 165.800 165.000 166.200 ;
        RECT 175.800 165.800 176.200 166.200 ;
        RECT 93.400 164.800 93.800 165.200 ;
        RECT 69.400 159.800 69.800 160.200 ;
        RECT 59.800 155.800 60.200 156.200 ;
        RECT 51.800 141.800 52.200 142.200 ;
        RECT 59.800 139.200 60.100 155.800 ;
        RECT 69.400 152.200 69.700 159.800 ;
        RECT 87.800 157.800 88.200 158.200 ;
        RECT 76.600 154.800 77.000 155.200 ;
        RECT 87.000 154.800 87.400 155.200 ;
        RECT 69.400 151.800 69.800 152.200 ;
        RECT 62.200 147.100 62.600 147.200 ;
        RECT 65.400 147.100 65.800 147.200 ;
        RECT 66.200 147.100 66.600 147.200 ;
        RECT 62.200 146.800 63.300 147.100 ;
        RECT 65.400 146.800 66.600 147.100 ;
        RECT 59.800 138.800 60.200 139.200 ;
        RECT 57.400 135.800 57.800 136.200 ;
        RECT 59.000 136.100 59.400 136.200 ;
        RECT 59.800 136.100 60.200 136.200 ;
        RECT 59.000 135.800 60.200 136.100 ;
        RECT 53.400 133.800 53.800 134.200 ;
        RECT 55.800 134.100 56.200 134.200 ;
        RECT 56.600 134.100 57.000 134.200 ;
        RECT 55.800 133.800 57.000 134.100 ;
        RECT 52.600 127.100 53.000 127.200 ;
        RECT 53.400 127.100 53.700 133.800 ;
        RECT 52.600 126.800 53.700 127.100 ;
        RECT 47.800 115.800 48.200 116.200 ;
        RECT 46.200 102.800 46.600 103.200 ;
        RECT 45.400 97.800 45.800 98.200 ;
        RECT 45.400 93.800 45.800 94.200 ;
        RECT 43.000 86.800 43.400 87.200 ;
        RECT 43.800 86.800 44.200 87.200 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 43.000 63.200 43.300 86.800 ;
        RECT 43.800 86.200 44.100 86.800 ;
        RECT 43.800 85.800 44.200 86.200 ;
        RECT 43.000 62.800 43.400 63.200 ;
        RECT 44.600 49.200 44.900 86.800 ;
        RECT 45.400 84.200 45.700 93.800 ;
        RECT 46.200 92.200 46.500 102.800 ;
        RECT 47.000 95.800 47.400 96.200 ;
        RECT 46.200 91.800 46.600 92.200 ;
        RECT 45.400 83.800 45.800 84.200 ;
        RECT 47.000 60.200 47.300 95.800 ;
        RECT 47.800 86.200 48.100 115.800 ;
        RECT 55.800 105.100 56.200 105.200 ;
        RECT 55.800 104.800 56.900 105.100 ;
        RECT 55.800 96.800 56.200 97.200 ;
        RECT 53.400 93.800 53.800 94.200 ;
        RECT 47.800 85.800 48.200 86.200 ;
        RECT 49.400 75.800 49.800 76.200 ;
        RECT 47.000 59.800 47.400 60.200 ;
        RECT 49.400 56.200 49.700 75.800 ;
        RECT 49.400 55.800 49.800 56.200 ;
        RECT 44.600 48.800 45.000 49.200 ;
        RECT 42.200 44.800 42.600 45.200 ;
        RECT 31.800 32.800 32.200 33.200 ;
        RECT 35.000 32.800 35.400 33.200 ;
        RECT 27.800 26.800 28.200 27.200 ;
        RECT 3.000 24.800 3.400 25.200 ;
        RECT 27.800 17.200 28.100 26.800 ;
        RECT 27.800 16.800 28.200 17.200 ;
        RECT 31.800 16.200 32.100 32.800 ;
        RECT 49.400 25.200 49.700 55.800 ;
        RECT 53.400 40.200 53.700 93.800 ;
        RECT 55.800 93.200 56.100 96.800 ;
        RECT 55.800 92.800 56.200 93.200 ;
        RECT 55.000 69.800 55.400 70.200 ;
        RECT 54.200 66.800 54.600 67.200 ;
        RECT 54.200 47.200 54.500 66.800 ;
        RECT 54.200 46.800 54.600 47.200 ;
        RECT 53.400 39.800 53.800 40.200 ;
        RECT 55.000 36.100 55.300 69.800 ;
        RECT 56.600 68.200 56.900 104.800 ;
        RECT 57.400 93.200 57.700 135.800 ;
        RECT 59.800 94.800 60.200 95.200 ;
        RECT 57.400 92.800 57.800 93.200 ;
        RECT 59.800 89.200 60.100 94.800 ;
        RECT 59.800 88.800 60.200 89.200 ;
        RECT 56.600 67.800 57.000 68.200 ;
        RECT 55.800 37.100 56.200 37.200 ;
        RECT 56.600 37.100 57.000 37.200 ;
        RECT 55.800 36.800 57.000 37.100 ;
        RECT 55.800 36.100 56.200 36.200 ;
        RECT 55.000 35.800 56.200 36.100 ;
        RECT 63.000 32.200 63.300 146.800 ;
        RECT 68.600 141.800 69.000 142.200 ;
        RECT 64.600 136.800 65.000 137.200 ;
        RECT 63.800 133.800 64.200 134.200 ;
        RECT 63.800 125.200 64.100 133.800 ;
        RECT 63.800 124.800 64.200 125.200 ;
        RECT 64.600 124.200 64.900 136.800 ;
        RECT 68.600 128.200 68.900 141.800 ;
        RECT 69.400 141.200 69.700 151.800 ;
        RECT 69.400 140.800 69.800 141.200 ;
        RECT 73.400 130.800 73.800 131.200 ;
        RECT 68.600 127.800 69.000 128.200 ;
        RECT 64.600 123.800 65.000 124.200 ;
        RECT 72.600 123.800 73.000 124.200 ;
        RECT 63.800 115.800 64.200 116.200 ;
        RECT 63.800 105.200 64.100 115.800 ;
        RECT 72.600 115.200 72.900 123.800 ;
        RECT 72.600 114.800 73.000 115.200 ;
        RECT 63.800 104.800 64.200 105.200 ;
        RECT 63.800 85.200 64.100 104.800 ;
        RECT 73.400 96.200 73.700 130.800 ;
        RECT 76.600 101.200 76.900 154.800 ;
        RECT 87.000 150.200 87.300 154.800 ;
        RECT 87.000 149.800 87.400 150.200 ;
        RECT 85.400 146.800 85.800 147.200 ;
        RECT 77.400 145.800 77.800 146.200 ;
        RECT 76.600 100.800 77.000 101.200 ;
        RECT 73.400 95.800 73.800 96.200 ;
        RECT 67.800 88.100 68.200 88.200 ;
        RECT 68.600 88.100 69.000 88.200 ;
        RECT 67.800 87.800 69.000 88.100 ;
        RECT 77.400 87.200 77.700 145.800 ;
        RECT 82.200 133.100 82.600 133.200 ;
        RECT 83.000 133.100 83.400 133.200 ;
        RECT 82.200 132.800 83.400 133.100 ;
        RECT 83.000 131.800 83.400 132.200 ;
        RECT 78.200 106.800 78.600 107.200 ;
        RECT 77.400 86.800 77.800 87.200 ;
        RECT 63.800 84.800 64.200 85.200 ;
        RECT 63.800 77.200 64.100 84.800 ;
        RECT 75.000 82.800 75.400 83.200 ;
        RECT 63.800 76.800 64.200 77.200 ;
        RECT 63.800 62.200 64.100 76.800 ;
        RECT 70.200 71.800 70.600 72.200 ;
        RECT 67.800 66.800 68.200 67.200 ;
        RECT 63.800 61.800 64.200 62.200 ;
        RECT 67.800 49.200 68.100 66.800 ;
        RECT 70.200 55.200 70.500 71.800 ;
        RECT 72.600 66.800 73.000 67.200 ;
        RECT 72.600 64.200 72.900 66.800 ;
        RECT 72.600 63.800 73.000 64.200 ;
        RECT 70.200 54.800 70.600 55.200 ;
        RECT 67.800 48.800 68.200 49.200 ;
        RECT 70.200 39.200 70.500 54.800 ;
        RECT 75.000 48.200 75.300 82.800 ;
        RECT 78.200 63.200 78.500 106.800 ;
        RECT 83.000 74.200 83.300 131.800 ;
        RECT 85.400 127.200 85.700 146.800 ;
        RECT 85.400 126.800 85.800 127.200 ;
        RECT 85.400 114.800 85.800 115.200 ;
        RECT 83.800 107.100 84.200 107.200 ;
        RECT 84.600 107.100 85.000 107.200 ;
        RECT 83.800 106.800 85.000 107.100 ;
        RECT 85.400 102.200 85.700 114.800 ;
        RECT 85.400 101.800 85.800 102.200 ;
        RECT 83.000 73.800 83.400 74.200 ;
        RECT 84.600 73.800 85.000 74.200 ;
        RECT 83.000 65.100 83.400 65.200 ;
        RECT 83.800 65.100 84.200 65.200 ;
        RECT 83.000 64.800 84.200 65.100 ;
        RECT 78.200 62.800 78.600 63.200 ;
        RECT 79.800 60.800 80.200 61.200 ;
        RECT 75.000 47.800 75.400 48.200 ;
        RECT 70.200 38.800 70.600 39.200 ;
        RECT 75.800 37.100 76.200 37.200 ;
        RECT 76.600 37.100 77.000 37.200 ;
        RECT 75.800 36.800 77.000 37.100 ;
        RECT 74.200 32.800 74.600 33.200 ;
        RECT 63.000 31.800 63.400 32.200 ;
        RECT 74.200 30.200 74.500 32.800 ;
        RECT 74.200 29.800 74.600 30.200 ;
        RECT 49.400 24.800 49.800 25.200 ;
        RECT 79.800 19.200 80.100 60.800 ;
        RECT 82.200 53.800 82.600 54.200 ;
        RECT 82.200 45.200 82.500 53.800 ;
        RECT 82.200 44.800 82.600 45.200 ;
        RECT 82.200 35.800 82.600 36.200 ;
        RECT 82.200 29.200 82.500 35.800 ;
        RECT 84.600 35.200 84.900 73.800 ;
        RECT 85.400 66.200 85.700 101.800 ;
        RECT 86.200 98.800 86.600 99.200 ;
        RECT 86.200 78.200 86.500 98.800 ;
        RECT 86.200 77.800 86.600 78.200 ;
        RECT 87.000 76.800 87.400 77.200 ;
        RECT 86.200 68.800 86.600 69.200 ;
        RECT 86.200 66.200 86.500 68.800 ;
        RECT 87.000 66.200 87.300 76.800 ;
        RECT 85.400 65.800 85.800 66.200 ;
        RECT 86.200 65.800 86.600 66.200 ;
        RECT 87.000 65.800 87.400 66.200 ;
        RECT 87.000 51.800 87.400 52.200 ;
        RECT 87.000 46.200 87.300 51.800 ;
        RECT 87.000 45.800 87.400 46.200 ;
        RECT 87.800 44.200 88.100 157.800 ;
        RECT 93.400 147.200 93.700 164.800 ;
        RECT 101.400 164.100 101.800 164.200 ;
        RECT 100.600 163.800 101.800 164.100 ;
        RECT 100.600 151.200 100.900 163.800 ;
        RECT 100.600 150.800 101.000 151.200 ;
        RECT 93.400 146.800 93.800 147.200 ;
        RECT 103.000 146.800 103.400 147.200 ;
        RECT 99.800 146.100 100.200 146.200 ;
        RECT 100.600 146.100 101.000 146.200 ;
        RECT 99.800 145.800 101.000 146.100 ;
        RECT 99.800 137.800 100.200 138.200 ;
        RECT 95.000 133.800 95.400 134.200 ;
        RECT 95.000 117.200 95.300 133.800 ;
        RECT 99.800 125.200 100.100 137.800 ;
        RECT 103.000 134.200 103.300 146.800 ;
        RECT 103.800 146.200 104.100 165.800 ;
        RECT 158.200 147.800 158.600 148.200 ;
        RECT 155.800 146.800 156.200 147.200 ;
        RECT 156.600 147.100 157.000 147.200 ;
        RECT 157.400 147.100 157.800 147.200 ;
        RECT 156.600 146.800 157.800 147.100 ;
        RECT 103.800 145.800 104.200 146.200 ;
        RECT 134.200 145.800 134.600 146.200 ;
        RECT 147.800 145.800 148.200 146.200 ;
        RECT 103.800 136.800 104.200 137.200 ;
        RECT 115.000 136.800 115.400 137.200 ;
        RECT 103.000 133.800 103.400 134.200 ;
        RECT 103.800 131.200 104.100 136.800 ;
        RECT 113.400 134.800 113.800 135.200 ;
        RECT 103.800 130.800 104.200 131.200 ;
        RECT 101.400 126.800 101.800 127.200 ;
        RECT 99.800 124.800 100.200 125.200 ;
        RECT 97.400 121.100 97.800 121.200 ;
        RECT 96.600 120.800 97.800 121.100 ;
        RECT 95.000 116.800 95.400 117.200 ;
        RECT 96.600 110.200 96.900 120.800 ;
        RECT 96.600 109.800 97.000 110.200 ;
        RECT 99.000 105.800 99.400 106.200 ;
        RECT 98.200 100.800 98.600 101.200 ;
        RECT 91.800 95.800 92.200 96.200 ;
        RECT 91.800 67.200 92.100 95.800 ;
        RECT 93.400 87.800 93.800 88.200 ;
        RECT 93.400 77.200 93.700 87.800 ;
        RECT 98.200 86.200 98.500 100.800 ;
        RECT 98.200 85.800 98.600 86.200 ;
        RECT 93.400 76.800 93.800 77.200 ;
        RECT 91.800 66.800 92.200 67.200 ;
        RECT 91.800 50.200 92.100 66.800 ;
        RECT 95.800 63.800 96.200 64.200 ;
        RECT 91.800 49.800 92.200 50.200 ;
        RECT 87.800 43.800 88.200 44.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 82.200 28.800 82.600 29.200 ;
        RECT 84.600 23.200 84.900 34.800 ;
        RECT 84.600 22.800 85.000 23.200 ;
        RECT 87.800 20.200 88.100 43.800 ;
        RECT 87.800 19.800 88.200 20.200 ;
        RECT 79.800 18.800 80.200 19.200 ;
        RECT 31.800 15.800 32.200 16.200 ;
        RECT 95.000 16.100 95.400 16.200 ;
        RECT 95.800 16.100 96.100 63.800 ;
        RECT 97.400 39.800 97.800 40.200 ;
        RECT 97.400 19.200 97.700 39.800 ;
        RECT 98.200 26.200 98.500 85.800 ;
        RECT 99.000 32.200 99.300 105.800 ;
        RECT 100.600 94.800 101.000 95.200 ;
        RECT 99.800 67.800 100.200 68.200 ;
        RECT 99.800 67.200 100.100 67.800 ;
        RECT 99.800 66.800 100.200 67.200 ;
        RECT 100.600 60.100 100.900 94.800 ;
        RECT 101.400 63.200 101.700 126.800 ;
        RECT 107.000 113.800 107.400 114.200 ;
        RECT 107.000 95.200 107.300 113.800 ;
        RECT 113.400 102.200 113.700 134.800 ;
        RECT 115.000 123.200 115.300 136.800 ;
        RECT 132.600 132.800 133.000 133.200 ;
        RECT 115.000 122.800 115.400 123.200 ;
        RECT 115.000 114.800 115.400 115.200 ;
        RECT 113.400 101.800 113.800 102.200 ;
        RECT 114.200 97.800 114.600 98.200 ;
        RECT 107.000 94.800 107.400 95.200 ;
        RECT 113.400 94.800 113.800 95.200 ;
        RECT 112.600 93.800 113.000 94.200 ;
        RECT 102.200 89.800 102.600 90.200 ;
        RECT 102.200 78.200 102.500 89.800 ;
        RECT 102.200 77.800 102.600 78.200 ;
        RECT 112.600 77.200 112.900 93.800 ;
        RECT 111.800 76.800 112.200 77.200 ;
        RECT 112.600 76.800 113.000 77.200 ;
        RECT 111.800 69.200 112.100 76.800 ;
        RECT 111.800 68.800 112.200 69.200 ;
        RECT 102.200 67.100 102.600 67.200 ;
        RECT 103.000 67.100 103.400 67.200 ;
        RECT 102.200 66.800 103.400 67.100 ;
        RECT 101.400 62.800 101.800 63.200 ;
        RECT 101.400 60.100 101.800 60.200 ;
        RECT 100.600 59.800 101.800 60.100 ;
        RECT 100.600 57.800 101.000 58.200 ;
        RECT 100.600 57.200 100.900 57.800 ;
        RECT 100.600 56.800 101.000 57.200 ;
        RECT 112.600 46.200 112.900 76.800 ;
        RECT 113.400 55.200 113.700 94.800 ;
        RECT 114.200 75.200 114.500 97.800 ;
        RECT 115.000 89.200 115.300 114.800 ;
        RECT 129.400 101.800 129.800 102.200 ;
        RECT 129.400 91.200 129.700 101.800 ;
        RECT 129.400 90.800 129.800 91.200 ;
        RECT 115.000 88.800 115.400 89.200 ;
        RECT 115.800 87.100 116.200 87.200 ;
        RECT 116.600 87.100 117.000 87.200 ;
        RECT 115.800 86.800 117.000 87.100 ;
        RECT 132.600 80.200 132.900 132.800 ;
        RECT 134.200 128.200 134.500 145.800 ;
        RECT 147.800 132.200 148.100 145.800 ;
        RECT 147.800 131.800 148.200 132.200 ;
        RECT 134.200 127.800 134.600 128.200 ;
        RECT 149.400 127.800 149.800 128.200 ;
        RECT 147.000 106.800 147.400 107.200 ;
        RECT 143.800 105.800 144.200 106.200 ;
        RECT 132.600 79.800 133.000 80.200 ;
        RECT 143.000 75.800 143.400 76.200 ;
        RECT 143.000 75.200 143.300 75.800 ;
        RECT 114.200 74.800 114.600 75.200 ;
        RECT 128.600 74.800 129.000 75.200 ;
        RECT 133.400 75.100 133.800 75.200 ;
        RECT 134.200 75.100 134.600 75.200 ;
        RECT 133.400 74.800 134.600 75.100 ;
        RECT 143.000 74.800 143.400 75.200 ;
        RECT 116.600 72.800 117.000 73.200 ;
        RECT 119.000 72.800 119.400 73.200 ;
        RECT 116.600 67.200 116.900 72.800 ;
        RECT 117.400 71.800 117.800 72.200 ;
        RECT 116.600 66.800 117.000 67.200 ;
        RECT 113.400 54.800 113.800 55.200 ;
        RECT 112.600 45.800 113.000 46.200 ;
        RECT 114.200 42.800 114.600 43.200 ;
        RECT 99.000 31.800 99.400 32.200 ;
        RECT 98.200 25.800 98.600 26.200 ;
        RECT 97.400 18.800 97.800 19.200 ;
        RECT 95.000 15.800 96.100 16.100 ;
        RECT 52.600 14.100 53.000 14.200 ;
        RECT 53.400 14.100 53.800 14.200 ;
        RECT 52.600 13.800 53.800 14.100 ;
        RECT 56.600 13.800 57.000 14.200 ;
        RECT 56.600 13.200 56.900 13.800 ;
        RECT 56.600 12.800 57.000 13.200 ;
        RECT 98.200 5.200 98.500 25.800 ;
        RECT 114.200 25.200 114.500 42.800 ;
        RECT 115.800 34.800 116.200 35.200 ;
        RECT 114.200 24.800 114.600 25.200 ;
        RECT 115.800 16.200 116.100 34.800 ;
        RECT 116.600 31.200 116.900 66.800 ;
        RECT 117.400 66.200 117.700 71.800 ;
        RECT 117.400 66.100 117.800 66.200 ;
        RECT 117.400 65.800 118.500 66.100 ;
        RECT 118.200 34.200 118.500 65.800 ;
        RECT 119.000 56.200 119.300 72.800 ;
        RECT 119.000 55.800 119.400 56.200 ;
        RECT 124.600 53.800 125.000 54.200 ;
        RECT 119.800 50.800 120.200 51.200 ;
        RECT 119.800 48.200 120.100 50.800 ;
        RECT 119.800 47.800 120.200 48.200 ;
        RECT 124.600 45.200 124.900 53.800 ;
        RECT 128.600 46.200 128.900 74.800 ;
        RECT 143.800 74.200 144.100 105.800 ;
        RECT 147.000 92.200 147.300 106.800 ;
        RECT 147.000 91.800 147.400 92.200 ;
        RECT 143.800 73.800 144.200 74.200 ;
        RECT 140.600 72.800 141.000 73.200 ;
        RECT 140.600 66.200 140.900 72.800 ;
        RECT 140.600 65.800 141.000 66.200 ;
        RECT 140.600 55.200 140.900 65.800 ;
        RECT 145.400 64.100 145.800 64.200 ;
        RECT 145.400 63.800 146.500 64.100 ;
        RECT 142.200 61.800 142.600 62.200 ;
        RECT 142.200 60.200 142.500 61.800 ;
        RECT 142.200 59.800 142.600 60.200 ;
        RECT 140.600 54.800 141.000 55.200 ;
        RECT 128.600 45.800 129.000 46.200 ;
        RECT 124.600 44.800 125.000 45.200 ;
        RECT 123.000 35.100 123.400 35.200 ;
        RECT 122.200 34.800 123.400 35.100 ;
        RECT 118.200 33.800 118.600 34.200 ;
        RECT 116.600 30.800 117.000 31.200 ;
        RECT 115.800 15.800 116.200 16.200 ;
        RECT 119.800 15.800 120.200 16.200 ;
        RECT 119.800 13.200 120.100 15.800 ;
        RECT 119.800 12.800 120.200 13.200 ;
        RECT 122.200 11.200 122.500 34.800 ;
        RECT 123.000 32.800 123.400 33.200 ;
        RECT 123.000 32.200 123.300 32.800 ;
        RECT 123.000 31.800 123.400 32.200 ;
        RECT 128.600 16.200 128.900 45.800 ;
        RECT 136.600 24.800 137.000 25.200 ;
        RECT 136.600 18.200 136.900 24.800 ;
        RECT 136.600 17.800 137.000 18.200 ;
        RECT 128.600 15.800 129.000 16.200 ;
        RECT 140.600 13.200 140.900 54.800 ;
        RECT 146.200 44.200 146.500 63.800 ;
        RECT 149.400 54.200 149.700 127.800 ;
        RECT 151.800 112.100 152.200 112.200 ;
        RECT 151.000 111.800 152.200 112.100 ;
        RECT 150.200 89.800 150.600 90.200 ;
        RECT 149.400 53.800 149.800 54.200 ;
        RECT 146.200 43.800 146.600 44.200 ;
        RECT 140.600 12.800 141.000 13.200 ;
        RECT 122.200 10.800 122.600 11.200 ;
        RECT 129.400 8.100 129.800 8.200 ;
        RECT 130.200 8.100 130.600 8.200 ;
        RECT 129.400 7.800 130.600 8.100 ;
        RECT 139.000 8.100 139.400 8.200 ;
        RECT 139.800 8.100 140.200 8.200 ;
        RECT 139.000 7.800 140.200 8.100 ;
        RECT 150.200 6.100 150.500 89.800 ;
        RECT 151.000 9.200 151.300 111.800 ;
        RECT 153.400 99.800 153.800 100.200 ;
        RECT 153.400 71.200 153.700 99.800 ;
        RECT 155.000 84.800 155.400 85.200 ;
        RECT 155.000 71.200 155.300 84.800 ;
        RECT 153.400 70.800 153.800 71.200 ;
        RECT 155.000 70.800 155.400 71.200 ;
        RECT 151.800 65.100 152.200 65.200 ;
        RECT 152.600 65.100 153.000 65.200 ;
        RECT 151.800 64.800 153.000 65.100 ;
        RECT 155.800 49.200 156.100 146.800 ;
        RECT 157.400 134.800 157.800 135.200 ;
        RECT 157.400 116.200 157.700 134.800 ;
        RECT 157.400 115.800 157.800 116.200 ;
        RECT 157.400 75.200 157.700 115.800 ;
        RECT 157.400 74.800 157.800 75.200 ;
        RECT 158.200 69.200 158.500 147.800 ;
        RECT 159.000 141.200 159.300 165.800 ;
        RECT 159.000 140.800 159.400 141.200 ;
        RECT 159.000 134.800 159.400 135.200 ;
        RECT 159.000 95.200 159.300 134.800 ;
        RECT 159.800 132.800 160.200 133.200 ;
        RECT 159.800 114.200 160.100 132.800 ;
        RECT 161.400 124.800 161.800 125.200 ;
        RECT 160.600 114.800 161.000 115.200 ;
        RECT 159.800 113.800 160.200 114.200 ;
        RECT 159.000 94.800 159.400 95.200 ;
        RECT 159.800 87.800 160.200 88.200 ;
        RECT 159.800 87.200 160.100 87.800 ;
        RECT 159.800 86.800 160.200 87.200 ;
        RECT 156.600 69.100 157.000 69.200 ;
        RECT 157.400 69.100 157.800 69.200 ;
        RECT 156.600 68.800 157.800 69.100 ;
        RECT 158.200 68.800 158.600 69.200 ;
        RECT 158.200 55.200 158.500 68.800 ;
        RECT 158.200 54.800 158.600 55.200 ;
        RECT 155.800 48.800 156.200 49.200 ;
        RECT 155.000 45.100 155.400 45.200 ;
        RECT 154.200 44.800 155.400 45.100 ;
        RECT 154.200 25.200 154.500 44.800 ;
        RECT 160.600 41.200 160.900 114.800 ;
        RECT 161.400 106.200 161.700 124.800 ;
        RECT 162.200 114.100 162.600 114.200 ;
        RECT 162.200 113.800 163.300 114.100 ;
        RECT 161.400 105.800 161.800 106.200 ;
        RECT 163.000 101.200 163.300 113.800 ;
        RECT 163.000 100.800 163.400 101.200 ;
        RECT 164.600 99.200 164.900 165.800 ;
        RECT 174.200 163.800 174.600 164.200 ;
        RECT 169.400 161.800 169.800 162.200 ;
        RECT 165.400 159.800 165.800 160.200 ;
        RECT 165.400 135.200 165.700 159.800 ;
        RECT 167.800 155.800 168.200 156.200 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 166.200 132.800 166.600 133.200 ;
        RECT 166.200 131.200 166.500 132.800 ;
        RECT 167.000 131.800 167.400 132.200 ;
        RECT 166.200 130.800 166.600 131.200 ;
        RECT 165.400 124.800 165.800 125.200 ;
        RECT 164.600 98.800 165.000 99.200 ;
        RECT 163.800 88.800 164.200 89.200 ;
        RECT 161.400 67.800 161.800 68.200 ;
        RECT 161.400 66.200 161.700 67.800 ;
        RECT 161.400 65.800 161.800 66.200 ;
        RECT 163.800 56.200 164.100 88.800 ;
        RECT 164.600 68.800 165.000 69.200 ;
        RECT 164.600 68.200 164.900 68.800 ;
        RECT 164.600 67.800 165.000 68.200 ;
        RECT 165.400 61.200 165.700 124.800 ;
        RECT 166.200 114.200 166.500 130.800 ;
        RECT 166.200 113.800 166.600 114.200 ;
        RECT 166.200 107.800 166.600 108.200 ;
        RECT 166.200 107.200 166.500 107.800 ;
        RECT 166.200 106.800 166.600 107.200 ;
        RECT 166.200 85.800 166.600 86.200 ;
        RECT 165.400 60.800 165.800 61.200 ;
        RECT 166.200 59.200 166.500 85.800 ;
        RECT 166.200 58.800 166.600 59.200 ;
        RECT 163.800 55.800 164.200 56.200 ;
        RECT 166.200 47.200 166.500 58.800 ;
        RECT 166.200 46.800 166.600 47.200 ;
        RECT 167.000 45.200 167.300 131.800 ;
        RECT 167.800 106.200 168.100 155.800 ;
        RECT 168.600 146.800 169.000 147.200 ;
        RECT 168.600 133.200 168.900 146.800 ;
        RECT 169.400 133.200 169.700 161.800 ;
        RECT 173.400 155.800 173.800 156.200 ;
        RECT 172.600 151.800 173.000 152.200 ;
        RECT 171.000 134.800 171.400 135.200 ;
        RECT 168.600 132.800 169.000 133.200 ;
        RECT 169.400 132.800 169.800 133.200 ;
        RECT 170.200 123.800 170.600 124.200 ;
        RECT 169.400 115.800 169.800 116.200 ;
        RECT 167.800 105.800 168.200 106.200 ;
        RECT 168.600 64.800 169.000 65.200 ;
        RECT 167.800 48.800 168.200 49.200 ;
        RECT 167.000 44.800 167.400 45.200 ;
        RECT 160.600 40.800 161.000 41.200 ;
        RECT 167.800 34.200 168.100 48.800 ;
        RECT 168.600 48.200 168.900 64.800 ;
        RECT 168.600 47.800 169.000 48.200 ;
        RECT 167.800 33.800 168.200 34.200 ;
        RECT 154.200 24.800 154.600 25.200 ;
        RECT 169.400 23.200 169.700 115.800 ;
        RECT 170.200 79.200 170.500 123.800 ;
        RECT 171.000 86.200 171.300 134.800 ;
        RECT 171.800 117.800 172.200 118.200 ;
        RECT 171.000 85.800 171.400 86.200 ;
        RECT 170.200 78.800 170.600 79.200 ;
        RECT 171.000 61.800 171.400 62.200 ;
        RECT 171.000 34.200 171.300 61.800 ;
        RECT 171.800 46.200 172.100 117.800 ;
        RECT 172.600 113.200 172.900 151.800 ;
        RECT 172.600 112.800 173.000 113.200 ;
        RECT 172.600 110.800 173.000 111.200 ;
        RECT 171.800 45.800 172.200 46.200 ;
        RECT 171.800 40.800 172.200 41.200 ;
        RECT 171.000 33.800 171.400 34.200 ;
        RECT 171.000 29.800 171.400 30.200 ;
        RECT 170.200 27.800 170.600 28.200 ;
        RECT 169.400 22.800 169.800 23.200 ;
        RECT 170.200 14.200 170.500 27.800 ;
        RECT 170.200 13.800 170.600 14.200 ;
        RECT 151.000 8.800 151.400 9.200 ;
        RECT 171.000 7.200 171.300 29.800 ;
        RECT 171.800 23.200 172.100 40.800 ;
        RECT 172.600 40.200 172.900 110.800 ;
        RECT 173.400 106.200 173.700 155.800 ;
        RECT 173.400 105.800 173.800 106.200 ;
        RECT 174.200 88.200 174.500 163.800 ;
        RECT 175.000 136.800 175.400 137.200 ;
        RECT 173.400 87.800 173.800 88.200 ;
        RECT 174.200 87.800 174.600 88.200 ;
        RECT 173.400 51.200 173.700 87.800 ;
        RECT 175.000 84.200 175.300 136.800 ;
        RECT 175.000 83.800 175.400 84.200 ;
        RECT 174.200 73.800 174.600 74.200 ;
        RECT 173.400 50.800 173.800 51.200 ;
        RECT 172.600 39.800 173.000 40.200 ;
        RECT 174.200 37.200 174.500 73.800 ;
        RECT 174.200 36.800 174.600 37.200 ;
        RECT 175.000 35.200 175.300 83.800 ;
        RECT 175.800 72.200 176.100 165.800 ;
        RECT 176.600 126.800 177.000 127.200 ;
        RECT 175.800 71.800 176.200 72.200 ;
        RECT 176.600 59.200 176.900 126.800 ;
        RECT 179.800 121.800 180.200 122.200 ;
        RECT 176.600 58.800 177.000 59.200 ;
        RECT 179.000 56.800 179.400 57.200 ;
        RECT 176.600 54.800 177.000 55.200 ;
        RECT 176.600 45.200 176.900 54.800 ;
        RECT 176.600 44.800 177.000 45.200 ;
        RECT 178.200 36.800 178.600 37.200 ;
        RECT 175.000 34.800 175.400 35.200 ;
        RECT 171.800 22.800 172.200 23.200 ;
        RECT 178.200 15.200 178.500 36.800 ;
        RECT 178.200 14.800 178.600 15.200 ;
        RECT 179.000 9.200 179.300 56.800 ;
        RECT 179.800 56.200 180.100 121.800 ;
        RECT 179.800 55.800 180.200 56.200 ;
        RECT 179.000 8.800 179.400 9.200 ;
        RECT 171.000 6.800 171.400 7.200 ;
        RECT 151.000 6.100 151.400 6.200 ;
        RECT 150.200 5.800 151.400 6.100 ;
        RECT 171.800 6.100 172.200 6.200 ;
        RECT 172.600 6.100 173.000 6.200 ;
        RECT 171.800 5.800 173.000 6.100 ;
        RECT 98.200 4.800 98.600 5.200 ;
      LAYER via4 ;
        RECT 24.600 85.800 25.000 86.200 ;
        RECT 42.200 132.800 42.600 133.200 ;
        RECT 49.400 146.800 49.800 147.200 ;
        RECT 66.200 146.800 66.600 147.200 ;
        RECT 56.600 36.800 57.000 37.200 ;
        RECT 68.600 87.800 69.000 88.200 ;
        RECT 84.600 106.800 85.000 107.200 ;
        RECT 83.800 64.800 84.200 65.200 ;
        RECT 134.200 74.800 134.600 75.200 ;
        RECT 152.600 64.800 153.000 65.200 ;
        RECT 157.400 68.800 157.800 69.200 ;
      LAYER metal5 ;
        RECT 45.400 147.100 45.800 147.200 ;
        RECT 49.400 147.100 49.800 147.200 ;
        RECT 45.400 146.800 49.800 147.100 ;
        RECT 66.200 147.100 66.600 147.200 ;
        RECT 156.600 147.100 157.000 147.200 ;
        RECT 66.200 146.800 157.000 147.100 ;
        RECT 99.800 146.100 100.200 146.200 ;
        RECT 100.500 146.100 101.000 146.200 ;
        RECT 99.800 145.800 101.000 146.100 ;
        RECT 100.500 145.700 101.000 145.800 ;
        RECT 31.000 136.100 31.400 136.200 ;
        RECT 59.000 136.100 59.400 136.200 ;
        RECT 31.000 135.800 59.400 136.100 ;
        RECT 34.200 134.100 34.600 134.200 ;
        RECT 55.800 134.100 56.200 134.200 ;
        RECT 34.200 133.800 56.200 134.100 ;
        RECT 42.200 133.100 42.600 133.200 ;
        RECT 82.200 133.100 82.600 133.200 ;
        RECT 42.200 132.800 82.600 133.100 ;
        RECT 172.600 112.800 173.000 113.200 ;
        RECT 172.600 112.200 172.900 112.800 ;
        RECT 172.500 111.700 173.000 112.200 ;
        RECT 84.600 107.100 85.000 107.200 ;
        RECT 166.200 107.100 166.600 107.200 ;
        RECT 84.600 106.800 166.600 107.100 ;
        RECT 68.600 88.100 69.000 88.200 ;
        RECT 159.800 88.100 160.200 88.200 ;
        RECT 68.600 87.800 160.200 88.100 ;
        RECT 43.800 87.100 44.200 87.200 ;
        RECT 115.800 87.100 116.200 87.200 ;
        RECT 43.800 86.800 116.200 87.100 ;
        RECT 24.600 86.100 25.000 86.200 ;
        RECT 33.400 86.100 33.800 86.200 ;
        RECT 24.600 85.800 33.800 86.100 ;
        RECT 134.200 75.100 134.600 75.200 ;
        RECT 143.000 75.100 143.400 75.200 ;
        RECT 134.200 74.800 143.400 75.100 ;
        RECT 157.400 69.100 157.800 69.200 ;
        RECT 164.600 69.100 165.000 69.200 ;
        RECT 157.400 68.800 165.000 69.100 ;
        RECT 99.800 67.800 100.200 68.200 ;
        RECT 99.800 67.100 100.100 67.800 ;
        RECT 102.200 67.100 102.600 67.200 ;
        RECT 99.800 66.800 102.600 67.100 ;
        RECT 83.800 65.100 84.200 65.200 ;
        RECT 152.600 65.100 153.000 65.200 ;
        RECT 83.800 64.800 153.000 65.100 ;
        RECT 100.500 58.700 101.000 59.200 ;
        RECT 100.600 58.200 100.900 58.700 ;
        RECT 100.600 57.800 101.000 58.200 ;
        RECT 56.600 37.100 57.000 37.200 ;
        RECT 75.800 37.100 76.200 37.200 ;
        RECT 56.600 36.800 76.200 37.100 ;
        RECT 74.200 33.100 74.600 33.200 ;
        RECT 74.200 32.800 123.300 33.100 ;
        RECT 123.000 32.200 123.300 32.800 ;
        RECT 123.000 31.800 123.400 32.200 ;
        RECT 52.600 14.100 53.000 14.200 ;
        RECT 56.600 14.100 57.000 14.200 ;
        RECT 52.600 13.800 57.000 14.100 ;
        RECT 129.400 8.100 129.800 8.200 ;
        RECT 139.000 8.100 139.400 8.200 ;
        RECT 129.400 7.800 139.400 8.100 ;
        RECT 171.800 6.100 172.200 6.200 ;
        RECT 172.500 6.100 173.000 6.200 ;
        RECT 171.800 5.800 173.000 6.100 ;
        RECT 172.500 5.700 173.000 5.800 ;
      LAYER metal6 ;
        RECT 100.500 58.700 101.000 146.200 ;
        RECT 172.500 5.700 173.000 112.200 ;
  END
END sram8t
END LIBRARY

