* NGSPICE file created from sram8t.ext - technology: scmos

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

.subckt sram8t vdd gnd clk rst_n cs re we addr[0] addr[1] addr[2] addr[3] din[0] din[1]
+ din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout[1] dout[2] dout[3] dout[4]
+ dout[5] dout[6] dout[7]
XMUX2X1_39 INVX1_49/Y INVX8_7/Y OR2X2_3/Y gnd MUX2X1_39/Y vdd MUX2X1
XMUX2X1_28 INVX1_59/Y INVX8_4/Y MUX2X1_29/S gnd MUX2X1_28/Y vdd MUX2X1
XMUX2X1_17 INVX1_18/Y INVX8_1/Y MUX2X1_10/S gnd MUX2X1_17/Y vdd MUX2X1
XNAND2X1_32 AOI22X1_10/Y NAND2X1_32/B gnd NOR3X1_11/C vdd NAND2X1
XNAND2X1_43 AOI22X1_15/Y NAND2X1_43/B gnd NOR3X1_15/C vdd NAND2X1
XNAND2X1_10 addr[3] INVX1_27/Y gnd INVX2_3/A vdd NAND2X1
XNAND2X1_54 INVX1_102/A NOR2X1_9/Y gnd NAND3X1_31/B vdd NAND2X1
XNAND2X1_21 AOI22X1_4/Y AOI22X1_5/Y gnd NOR3X1_7/C vdd NAND2X1
XOAI22X1_3 INVX1_33/Y INVX4_5/Y OAI22X1_4/C INVX1_34/Y gnd NOR3X1_8/C vdd OAI22X1
XFILL_11_1_0 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XDFFPOSX1_125 NOR2X1_24/A CLKBUF1_2/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_103 INVX1_63/A CLKBUF1_1/Y MUX2X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 NOR2X1_30/A CLKBUF1_9/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XFILL_0_0_0 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XMUX2X1_29 INVX1_60/Y INVX8_5/Y MUX2X1_29/S gnd MUX2X1_29/Y vdd MUX2X1
XMUX2X1_18 INVX8_6/Y INVX1_40/Y MUX2X1_18/S gnd MUX2X1_18/Y vdd MUX2X1
XNAND2X1_44 NOR2X1_43/A AND2X2_2/A gnd NAND3X1_23/A vdd NAND2X1
XNAND2X1_33 NOR2X1_32/A INVX2_5/A gnd NAND3X1_15/B vdd NAND2X1
XNAND2X1_11 INVX1_26/Y INVX2_3/Y gnd OR2X2_3/A vdd NAND2X1
XNAND2X1_55 AOI22X1_22/Y NAND2X1_55/B gnd NOR3X1_19/C vdd NAND2X1
XAOI22X1_1 INVX1_43/A INVX1_105/A INVX1_79/A NOR2X1_8/Y gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_22 NOR2X1_30/A INVX2_5/A gnd NAND3X1_8/B vdd NAND2X1
XAOI22X1_20 NOR2X1_26/A AND2X2_1/A NOR2X1_1/Y INVX1_17/A gnd AOI22X1_20/Y vdd AOI22X1
XOAI22X1_4 INVX1_37/Y INVX4_5/Y OAI22X1_4/C INVX1_38/Y gnd OAI22X1_4/Y vdd OAI22X1
XFILL_11_1_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XDFFPOSX1_115 NOR2X1_31/A CLKBUF1_4/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_104 INVX1_64/A CLKBUF1_9/Y MUX2X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_126 NOR2X1_25/A CLKBUF1_3/Y AOI21X1_14/Y gnd vdd DFFPOSX1
XFILL_10_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XAOI22X1_2 NOR2X1_9/Y INVX1_95/A INVX1_65/A INVX1_45/A gnd AOI22X1_2/Y vdd AOI22X1
XNAND2X1_23 INVX1_59/A NOR2X1_5/Y gnd OAI21X1_6/C vdd NAND2X1
XMUX2X1_19 INVX8_1/Y INVX1_54/Y MUX2X1_18/S gnd MUX2X1_19/Y vdd MUX2X1
XNAND2X1_34 INVX1_83/A NOR2X1_8/Y gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_12 INVX1_57/A NOR2X1_5/Y gnd OAI21X1_2/C vdd NAND2X1
XNAND2X1_45 NOR2X1_33/A INVX2_5/A gnd NAND2X1_45/Y vdd NAND2X1
XNAND2X1_56 INVX4_1/Y NOR2X1_5/Y gnd MUX2X1_29/S vdd NAND2X1
XAOI22X1_21 NOR2X1_37/A INVX4_5/A NOR2X1_5/Y INVX1_64/A gnd NAND3X1_31/C vdd AOI22X1
XAOI22X1_10 INVX1_43/A INVX1_108/A INVX1_82/A NOR2X1_8/Y gnd AOI22X1_10/Y vdd AOI22X1
XOAI22X1_5 INVX1_41/Y OR2X2_3/A INVX1_43/Y INVX1_42/Y gnd NOR3X1_12/C vdd OAI22X1
XDFFPOSX1_105 INVX1_21/A DFFSR_1/CLK MUX2X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_116 NOR2X1_32/A CLKBUF1_9/Y AOI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_127 NOR2X1_26/A CLKBUF1_10/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XINVX8_1 din[7] gnd INVX8_1/Y vdd INVX8
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XAOI22X1_3 NOR2X1_20/A AND2X2_1/A NOR2X1_1/Y INVX1_11/A gnd AOI22X1_3/Y vdd AOI22X1
XAOI22X1_11 NOR2X1_9/Y INVX1_98/A INVX1_68/A INVX1_45/A gnd NAND2X1_32/B vdd AOI22X1
XNAND2X1_13 INVX1_71/A NOR2X1_6/Y gnd NAND3X1_3/B vdd NAND2X1
XNAND2X1_24 INVX1_73/A NOR2X1_6/Y gnd NAND2X1_24/Y vdd NAND2X1
XNAND2X1_57 INVX4_1/Y INVX1_45/A gnd MUX2X1_45/S vdd NAND2X1
XNAND2X1_46 INVX1_63/A NOR2X1_5/Y gnd NAND2X1_46/Y vdd NAND2X1
XAOI22X1_22 NOR2X1_27/A AND2X2_1/A NOR2X1_6/Y INVX1_78/A gnd AOI22X1_22/Y vdd AOI22X1
XNOR3X1_1 addr[0] INVX1_2/Y INVX4_2/A gnd INVX1_43/A vdd NOR3X1
XNAND2X1_35 INVX1_75/A NOR2X1_6/Y gnd NAND2X1_35/Y vdd NAND2X1
XFILL_6_2_0 gnd vdd FILL
XOAI22X1_6 INVX1_47/Y INVX4_5/Y OAI22X1_4/C INVX1_48/Y gnd OAI22X1_6/Y vdd OAI22X1
XFILL_14_1_0 gnd vdd FILL
XDFFPOSX1_106 INVX1_29/A CLKBUF1_4/Y MUX2X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_117 INVX1_40/A CLKBUF1_4/Y MUX2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 NOR2X1_27/A CLKBUF1_10/Y AOI21X1_16/Y gnd vdd DFFPOSX1
XINVX8_2 din[0] gnd INVX8_2/Y vdd INVX8
XFILL_3_0_0 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XAOI22X1_4 INVX1_43/A INVX1_106/A INVX1_80/A NOR2X1_8/Y gnd AOI22X1_4/Y vdd AOI22X1
XNAND2X1_25 INVX1_89/A NOR2X1_7/Y gnd NAND3X1_10/C vdd NAND2X1
XNAND2X1_47 NOR2X1_44/A AND2X2_2/A gnd NAND3X1_25/A vdd NAND2X1
XNAND2X1_14 INVX1_87/A NOR2X1_7/Y gnd NAND3X1_3/C vdd NAND2X1
XAOI22X1_12 NOR2X1_23/A AND2X2_1/A NOR2X1_1/Y INVX1_14/A gnd AOI22X1_12/Y vdd AOI22X1
XNOR3X1_2 NOR3X1_2/A addr[1] NOR2X1_5/A gnd INVX4_5/A vdd NOR3X1
XAOI22X1_23 INVX1_104/A INVX4_4/A NOR2X1_7/Y INVX1_94/A gnd NAND2X1_55/B vdd AOI22X1
XNAND2X1_58 INVX4_1/Y NOR2X1_6/Y gnd MUX2X1_52/S vdd NAND2X1
XNAND2X1_36 INVX1_15/A NOR2X1_1/Y gnd NAND2X1_36/Y vdd NAND2X1
XOAI22X1_7 INVX1_51/Y INVX4_5/Y OAI22X1_4/C INVX1_52/Y gnd NOR3X1_16/C vdd OAI22X1
XFILL_14_1_1 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XDFFPOSX1_107 INVX1_33/A DFFSR_1/CLK MUX2X1_22/Y gnd vdd DFFPOSX1
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_118 NOR2X1_33/A CLKBUF1_3/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XINVX8_3 din[1] gnd INVX8_3/Y vdd INVX8
XFILL_3_0_1 gnd vdd FILL
XNAND2X1_48 INVX1_93/A NOR2X1_7/Y gnd NAND3X1_25/C vdd NAND2X1
XNAND2X1_26 AOI22X1_7/Y AOI22X1_8/Y gnd NOR3X1_9/C vdd NAND2X1
XNAND2X1_15 AOI22X1_1/Y AOI22X1_2/Y gnd NOR3X1_5/C vdd NAND2X1
XAOI22X1_13 NOR2X1_36/A INVX4_5/A NOR2X1_5/Y INVX1_61/A gnd NAND3X1_19/C vdd AOI22X1
XNAND2X1_37 INVX1_99/A NOR2X1_9/Y gnd NAND3X1_19/B vdd NAND2X1
XAOI22X1_5 NOR2X1_9/Y INVX1_96/A INVX1_66/A INVX1_45/A gnd AOI22X1_5/Y vdd AOI22X1
XNAND2X1_59 INVX4_1/Y NOR2X1_8/Y gnd MUX2X1_70/S vdd NAND2X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XOAI22X1_8 INVX1_55/Y OR2X2_3/A INVX1_43/Y INVX1_1/Y gnd NOR3X1_18/C vdd OAI22X1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XDFFPOSX1_108 INVX1_37/A DFFSR_1/CLK MUX2X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_119 NOR2X1_34/A CLKBUF1_10/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XMUX2X1_1 INVX1_1/Y INVX8_1/Y MUX2X1_1/S gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_90 NOR2X1_39/A CLKBUF1_8/Y AOI21X1_26/Y gnd vdd DFFPOSX1
XINVX8_4 din[2] gnd INVX8_4/Y vdd INVX8
XFILL_12_2_0 gnd vdd FILL
XNAND3X1_1 INVX4_2/Y INVX4_1/Y INVX4_3/Y gnd MUX2X1_2/S vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XNAND2X1_27 NOR2X1_40/A AND2X2_2/A gnd NAND3X1_11/A vdd NAND2X1
XNAND2X1_49 AOI22X1_18/Y AOI22X1_19/Y gnd NOR3X1_17/C vdd NAND2X1
XNAND2X1_16 NOR2X1_38/A AND2X2_2/A gnd NAND3X1_4/A vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XAOI22X1_6 AOI22X1_6/A AND2X2_1/A NOR2X1_1/Y INVX1_12/A gnd AOI22X1_6/Y vdd AOI22X1
XNAND2X1_38 INVX1_103/A INVX4_4/A gnd NAND2X1_38/Y vdd NAND2X1
XAOI22X1_14 NOR2X1_24/A AND2X2_1/A AND2X2_2/A NOR2X1_42/A gnd NAND3X1_20/A vdd AOI22X1
XNOR3X1_4 NOR3X1_4/A addr[2] INVX2_1/A gnd AND2X2_2/A vdd NOR3X1
XMUX2X1_2 INVX1_3/Y INVX8_2/Y MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XDFFPOSX1_109 NOR2X1_36/A CLKBUF1_5/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XFILL_6_0_0 gnd vdd FILL
XDFFPOSX1_91 NOR2X1_40/A CLKBUF1_8/Y AOI21X1_27/Y gnd vdd DFFPOSX1
XINVX8_5 din[3] gnd INVX8_5/Y vdd INVX8
XDFFPOSX1_80 INVX1_56/A CLKBUF1_9/Y MUX2X1_49/Y gnd vdd DFFPOSX1
XFILL_12_2_1 gnd vdd FILL
XNAND3X1_2 INVX1_3/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_3/A vdd NAND3X1
XNAND2X1_28 NOR2X1_31/A INVX2_5/A gnd NAND2X1_28/Y vdd NAND2X1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_17 NOR2X1_29/A INVX2_5/A gnd NAND3X1_4/B vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XAOI22X1_7 INVX1_43/A AOI22X1_7/B INVX1_81/A NOR2X1_8/Y gnd AOI22X1_7/Y vdd AOI22X1
XNAND2X1_39 INVX1_91/A NOR2X1_7/Y gnd NAND2X1_39/Y vdd NAND2X1
XNOR3X1_5 NOR3X1_5/A NOR3X1_5/B NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XAOI22X1_15 INVX1_43/A INVX1_109/A INVX1_84/A NOR2X1_8/Y gnd AOI22X1_15/Y vdd AOI22X1
XMUX2X1_3 INVX1_4/Y INVX8_3/Y MUX2X1_2/S gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XDFFPOSX1_70 INVX1_76/A CLKBUF1_8/Y MUX2X1_55/Y gnd vdd DFFPOSX1
XDFFPOSX1_92 NOR2X1_41/A CLKBUF1_2/Y AOI21X1_28/Y gnd vdd DFFPOSX1
XINVX8_6 din[4] gnd INVX8_6/Y vdd INVX8
XDFFPOSX1_81 INVX1_25/A DFFSR_8/CLK MUX2X1_34/Y gnd vdd DFFPOSX1
XAOI22X1_8 NOR2X1_9/Y INVX1_97/A INVX1_67/A INVX1_45/A gnd AOI22X1_8/Y vdd AOI22X1
XNAND3X1_3 NAND3X1_3/A NAND3X1_3/B NAND3X1_3/C gnd NOR3X1_5/A vdd NAND3X1
XAOI22X1_16 NOR2X1_9/Y INVX1_100/A INVX1_69/A INVX1_45/A gnd NAND2X1_43/B vdd AOI22X1
XNAND2X1_29 INVX1_60/A NOR2X1_5/Y gnd OAI21X1_8/C vdd NAND2X1
XNOR3X1_6 NOR3X1_6/A NOR3X1_6/B NOR3X1_6/C gnd NOR3X1_6/Y vdd NOR3X1
XNAND2X1_18 INVX1_58/A NOR2X1_5/Y gnd OAI21X1_4/C vdd NAND2X1
XMUX2X1_4 INVX1_5/Y INVX8_4/Y MUX2X1_2/S gnd MUX2X1_4/Y vdd MUX2X1
XFILL_17_1 gnd vdd FILL
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XDFFPOSX1_60 INVX1_38/A CLKBUF1_5/Y MUX2X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_93 NOR2X1_42/A CLKBUF1_3/Y AOI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_82 INVX1_31/A CLKBUF1_1/Y MUX2X1_35/Y gnd vdd DFFPOSX1
XINVX8_7 din[5] gnd INVX8_7/Y vdd INVX8
XDFFPOSX1_71 INVX1_77/A CLKBUF1_10/Y MUX2X1_56/Y gnd vdd DFFPOSX1
XFILL_15_2_0 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XAOI22X1_9 AOI22X1_9/A AND2X2_1/A NOR2X1_1/Y INVX1_13/A gnd AOI22X1_9/Y vdd AOI22X1
XNAND3X1_4 NAND3X1_4/A NAND3X1_4/B AOI22X1_3/Y gnd NOR3X1_5/B vdd NAND3X1
XNAND2X1_19 NOR2X1_39/A AND2X2_2/A gnd NAND3X1_6/A vdd NAND2X1
XNOR3X1_7 NOR3X1_7/A NOR3X1_7/B NOR3X1_7/C gnd NOR3X1_7/Y vdd NOR3X1
XAOI22X1_17 NOR2X1_25/A AND2X2_1/A NOR2X1_1/Y INVX1_16/A gnd AOI22X1_17/Y vdd AOI22X1
XOAI21X1_1 INVX4_4/Y INVX1_20/Y NOR2X1_3/B gnd NOR3X1_3/B vdd OAI21X1
XFILL_9_0_0 gnd vdd FILL
XMUX2X1_5 INVX1_6/Y INVX8_5/Y MUX2X1_2/S gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 clk gnd DFFSR_8/CLK vdd CLKBUF1
XINVX8_8 din[6] gnd INVX8_8/Y vdd INVX8
XFILL_15_2_1 gnd vdd FILL
XDFFPOSX1_94 NOR2X1_43/A CLKBUF1_8/Y AOI21X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_72 INVX1_78/A CLKBUF1_10/Y MUX2X1_57/Y gnd vdd DFFPOSX1
XDFFPOSX1_83 INVX1_35/A DFFSR_8/CLK MUX2X1_36/Y gnd vdd DFFPOSX1
XDFFPOSX1_50 INVX1_80/A CLKBUF1_9/Y MUX2X1_65/Y gnd vdd DFFPOSX1
XDFFPOSX1_61 NOR2X1_47/A CLKBUF1_9/Y AOI21X1_33/Y gnd vdd DFFPOSX1
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XNAND3X1_5 INVX1_4/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_5/Y vdd NAND3X1
XAOI22X1_18 INVX1_43/A INVX1_110/A INVX1_85/A NOR2X1_8/Y gnd AOI22X1_18/Y vdd AOI22X1
XNOR3X1_8 NOR3X1_8/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XFILL_9_0_1 gnd vdd FILL
XOAI21X1_2 OR2X2_3/A INVX1_25/Y OAI21X1_2/C gnd NOR3X1_3/A vdd OAI21X1
XMUX2X1_6 INVX1_7/Y INVX8_6/Y MUX2X1_2/S gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 clk gnd CLKBUF1_7/Y vdd CLKBUF1
XDFFPOSX1_73 INVX1_65/A CLKBUF1_5/Y MUX2X1_42/Y gnd vdd DFFPOSX1
XDFFPOSX1_95 NOR2X1_44/A CLKBUF1_8/Y AOI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_84 INVX1_39/A DFFSR_1/CLK MUX2X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_62 INVX1_48/A CLKBUF1_4/Y MUX2X1_62/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 INVX1_81/A CLKBUF1_9/Y MUX2X1_66/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 INVX1_102/A CLKBUF1_7/Y MUX2X1_87/Y gnd vdd DFFPOSX1
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XNAND3X1_6 NAND3X1_6/A NAND3X1_5/Y NAND3X1_6/C gnd NOR3X1_7/A vdd NAND3X1
XNOR3X1_9 NOR3X1_9/A NOR3X1_9/B NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XAOI22X1_19 NOR2X1_9/Y INVX1_101/A INVX1_70/A INVX1_45/A gnd AOI22X1_19/Y vdd AOI22X1
XAOI21X1_30 INVX8_7/Y AND2X2_2/Y NOR2X1_43/Y gnd AOI21X1_30/Y vdd AOI21X1
XOAI21X1_3 INVX4_4/Y INVX1_28/Y NOR2X1_3/B gnd NOR3X1_6/B vdd OAI21X1
XMUX2X1_7 INVX1_8/Y INVX8_7/Y MUX2X1_2/S gnd MUX2X1_7/Y vdd MUX2X1
XCLKBUF1_8 clk gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XDFFPOSX1_41 INVX1_87/A CLKBUF1_2/Y MUX2X1_72/Y gnd vdd DFFPOSX1
XDFFPOSX1_52 INVX1_82/A CLKBUF1_9/Y MUX2X1_67/Y gnd vdd DFFPOSX1
XDFFPOSX1_63 INVX1_52/A DFFSR_8/CLK MUX2X1_63/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 INVX1_46/A DFFSR_8/CLK MUX2X1_93/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 INVX1_66/A CLKBUF1_7/Y MUX2X1_43/Y gnd vdd DFFPOSX1
XDFFPOSX1_85 INVX1_41/A DFFSR_8/CLK MUX2X1_38/Y gnd vdd DFFPOSX1
XDFFPOSX1_96 NOR2X1_45/A CLKBUF1_3/Y AOI21X1_32/Y gnd vdd DFFPOSX1
XFILL_15_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XNAND3X1_7 INVX1_72/A INVX2_4/Y INVX2_3/Y gnd NAND3X1_7/Y vdd NAND3X1
XBUFX2_1 DFFSR_1/Q gnd dout[0] vdd BUFX2
XAOI21X1_1 NOR3X1_3/Y NOR3X1_5/Y NOR2X1_3/Y gnd DFFSR_1/D vdd AOI21X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_31 INVX8_8/Y AND2X2_2/Y NOR2X1_44/Y gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_20 INVX8_5/Y MUX2X1_18/S NOR2X1_32/Y gnd AOI21X1_20/Y vdd AOI21X1
XOAI21X1_4 OR2X2_3/A INVX1_31/Y OAI21X1_4/C gnd NOR3X1_6/A vdd OAI21X1
XMUX2X1_8 INVX1_9/Y INVX8_8/Y MUX2X1_2/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XCLKBUF1_9 clk gnd CLKBUF1_9/Y vdd CLKBUF1
XDFFPOSX1_42 INVX1_88/A CLKBUF1_5/Y MUX2X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 INVX1_67/A CLKBUF1_5/Y MUX2X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_64 NOR2X1_48/A CLKBUF1_7/Y AOI21X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 INVX1_49/A CLKBUF1_1/Y MUX2X1_39/Y gnd vdd DFFPOSX1
XDFFPOSX1_53 INVX1_83/A CLKBUF1_1/Y MUX2X1_68/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 INVX1_108/A CLKBUF1_9/Y MUX2X1_99/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 INVX1_50/A DFFSR_8/CLK MUX2X1_94/Y gnd vdd DFFPOSX1
XDFFPOSX1_97 INVX1_57/A DFFSR_8/CLK MUX2X1_26/Y gnd vdd DFFPOSX1
XFILL_15_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XBUFX2_2 BUFX2_2/A gnd dout[1] vdd BUFX2
XNAND3X1_8 NAND3X1_7/Y NAND3X1_8/B AOI22X1_6/Y gnd NOR3X1_7/B vdd NAND3X1
XAOI21X1_2 NOR3X1_6/Y NOR3X1_7/Y AOI21X1_2/C gnd DFFSR_2/D vdd AOI21X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XOAI21X1_5 INVX4_4/Y INVX1_32/Y NOR2X1_3/B gnd NOR3X1_8/B vdd OAI21X1
XAOI21X1_10 INVX8_3/Y AND2X2_1/Y NOR2X1_21/Y gnd AOI21X1_10/Y vdd AOI21X1
XAOI21X1_21 INVX8_7/Y MUX2X1_18/S NOR2X1_33/Y gnd AOI21X1_21/Y vdd AOI21X1
XAOI21X1_32 INVX8_1/Y AND2X2_2/Y NOR2X1_45/Y gnd AOI21X1_32/Y vdd AOI21X1
XMUX2X1_9 INVX1_10/Y INVX8_1/Y MUX2X1_2/S gnd MUX2X1_9/Y vdd MUX2X1
XDFFPOSX1_76 INVX1_68/A CLKBUF1_5/Y MUX2X1_45/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 INVX1_89/A CLKBUF1_2/Y MUX2X1_74/Y gnd vdd DFFPOSX1
XDFFPOSX1_65 INVX1_71/A CLKBUF1_8/Y MUX2X1_50/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 INVX1_4/A CLKBUF1_2/Y MUX2X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_54 INVX1_84/A CLKBUF1_7/Y MUX2X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_87 INVX1_53/A CLKBUF1_1/Y MUX2X1_40/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX1_58/A CLKBUF1_1/Y MUX2X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_32 INVX1_104/A CLKBUF1_10/Y MUX2X1_95/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 INVX1_42/A CLKBUF1_7/Y MUX2X1_100/Y gnd vdd DFFPOSX1
XNOR3X1_10 OAI21X1_8/Y NOR3X1_10/B OAI22X1_4/Y gnd AOI21X1_4/A vdd NOR3X1
XBUFX2_3 DFFSR_3/Q gnd dout[2] vdd BUFX2
XNAND3X1_9 INVX1_5/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_9/Y vdd NAND3X1
XAOI21X1_3 NOR3X1_8/Y NOR3X1_9/Y AOI21X1_3/C gnd DFFSR_3/D vdd AOI21X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XNOR2X1_1 INVX4_2/A OR2X2_2/Y gnd NOR2X1_1/Y vdd NOR2X1
XAOI21X1_11 INVX8_4/Y AND2X2_1/Y NOR2X1_22/Y gnd AOI21X1_11/Y vdd AOI21X1
XAOI21X1_22 INVX8_8/Y MUX2X1_18/S NOR2X1_34/Y gnd AOI21X1_22/Y vdd AOI21X1
XOAI21X1_6 OR2X2_3/A INVX1_35/Y OAI21X1_6/C gnd NOR3X1_8/A vdd OAI21X1
XAOI21X1_33 INVX8_6/Y NOR2X1_48/B NOR2X1_47/Y gnd AOI21X1_33/Y vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XDFFPOSX1_11 INVX1_5/A CLKBUF1_2/Y MUX2X1_4/Y gnd vdd DFFPOSX1
XDFFPOSX1_33 INVX1_95/A CLKBUF1_5/Y MUX2X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 INVX1_90/A CLKBUF1_2/Y MUX2X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 INVX1_55/A CLKBUF1_4/Y MUX2X1_41/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 INVX1_85/A CLKBUF1_4/Y MUX2X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 INVX1_109/A CLKBUF1_7/Y MUX2X1_101/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_66 INVX1_72/A CLKBUF1_10/Y MUX2X1_51/Y gnd vdd DFFPOSX1
XDFFPOSX1_99 INVX1_59/A CLKBUF1_1/Y MUX2X1_28/Y gnd vdd DFFPOSX1
XDFFPOSX1_77 INVX1_44/A CLKBUF1_1/Y MUX2X1_46/Y gnd vdd DFFPOSX1
XNOR3X1_11 NOR3X1_11/A NOR3X1_11/B NOR3X1_11/C gnd NOR3X1_11/Y vdd NOR3X1
XBUFX2_4 BUFX2_4/A gnd dout[3] vdd BUFX2
XAOI21X1_4 AOI21X1_4/A NOR3X1_11/Y AOI21X1_4/C gnd DFFSR_4/D vdd AOI21X1
XINVX2_4 OR2X2_2/Y gnd INVX2_4/Y vdd INVX2
XNOR2X1_2 we NOR2X1_2/B gnd NOR2X1_3/B vdd NOR2X1
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XOAI21X1_7 INVX4_4/Y INVX1_36/Y NOR2X1_3/B gnd NOR3X1_10/B vdd OAI21X1
XAOI21X1_23 INVX8_6/Y MUX2X1_20/S NOR2X1_36/Y gnd AOI21X1_23/Y vdd AOI21X1
XAOI21X1_12 INVX8_5/Y AND2X2_1/Y NOR2X1_23/Y gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_34 INVX8_1/Y NOR2X1_48/B NOR2X1_48/Y gnd AOI21X1_34/Y vdd AOI21X1
XFILL_13_1_1 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_78 INVX1_69/A CLKBUF1_5/Y MUX2X1_47/Y gnd vdd DFFPOSX1
XDFFPOSX1_67 INVX1_73/A CLKBUF1_8/Y MUX2X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_12 INVX1_6/A CLKBUF1_2/Y MUX2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_89 NOR2X1_38/A CLKBUF1_2/Y AOI21X1_25/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XDFFPOSX1_56 INVX1_86/A CLKBUF1_1/Y MUX2X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 INVX1_110/A CLKBUF1_9/Y MUX2X1_102/Y gnd vdd DFFPOSX1
XDFFPOSX1_45 INVX1_91/A CLKBUF1_3/Y MUX2X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_34 INVX1_96/A CLKBUF1_7/Y MUX2X1_81/Y gnd vdd DFFPOSX1
XNOR3X1_12 NOR3X1_12/A OAI21X1_9/Y NOR3X1_12/C gnd NOR3X1_12/Y vdd NOR3X1
XBUFX2_5 BUFX2_5/A gnd dout[4] vdd BUFX2
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XAOI21X1_5 NOR3X1_12/Y NOR3X1_13/Y AOI21X1_5/C gnd DFFSR_5/D vdd AOI21X1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XNOR2X1_3 DFFSR_1/Q NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_13 INVX8_6/Y AND2X2_1/Y NOR2X1_24/Y gnd AOI21X1_13/Y vdd AOI21X1
XAOI21X1_24 INVX8_1/Y MUX2X1_20/S NOR2X1_37/Y gnd AOI21X1_24/Y vdd AOI21X1
XOAI21X1_8 OR2X2_3/A INVX1_39/Y OAI21X1_8/C gnd OAI21X1_8/Y vdd OAI21X1
XDFFPOSX1_46 INVX1_92/A CLKBUF1_8/Y MUX2X1_77/Y gnd vdd DFFPOSX1
XDFFPOSX1_57 INVX1_22/A DFFSR_1/CLK MUX2X1_58/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 INVX1_7/A CLKBUF1_2/Y MUX2X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 INVX1_97/A CLKBUF1_5/Y MUX2X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_79 INVX1_70/A CLKBUF1_4/Y MUX2X1_48/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 INVX1_74/A CLKBUF1_10/Y MUX2X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 INVX1_1/A CLKBUF1_7/Y MUX2X1_1/Y gnd vdd DFFPOSX1
XFILL_11_2_0 gnd vdd FILL
XNOR3X1_13 NOR3X1_13/A NOR3X1_13/B NOR3X1_13/C gnd NOR3X1_13/Y vdd NOR3X1
XBUFX2_6 BUFX2_6/A gnd dout[5] vdd BUFX2
XNAND2X1_1 we cs gnd INVX4_1/A vdd NAND2X1
XFILL_16_1_0 gnd vdd FILL
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XDFFPOSX1_1 INVX1_11/A CLKBUF1_2/Y MUX2X1_10/Y gnd vdd DFFPOSX1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XFILL_8_2_0 gnd vdd FILL
XAOI21X1_6 NOR3X1_14/Y AOI21X1_6/B AOI21X1_6/C gnd DFFSR_6/D vdd AOI21X1
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_4 INVX2_1/A INVX4_2/A gnd INVX4_4/A vdd NOR2X1
XAOI21X1_25 INVX8_2/Y AND2X2_2/Y NOR2X1_38/Y gnd AOI21X1_25/Y vdd AOI21X1
XAOI21X1_14 INVX8_7/Y AND2X2_1/Y NOR2X1_25/Y gnd AOI21X1_14/Y vdd AOI21X1
XOAI21X1_9 INVX2_5/Y INVX1_40/Y NOR2X1_3/B gnd OAI21X1_9/Y vdd OAI21X1
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_36 INVX1_98/A CLKBUF1_5/Y MUX2X1_83/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 INVX1_8/A CLKBUF1_8/Y MUX2X1_7/Y gnd vdd DFFPOSX1
XDFFPOSX1_47 INVX1_93/A CLKBUF1_8/Y MUX2X1_78/Y gnd vdd DFFPOSX1
XDFFPOSX1_25 INVX1_20/A DFFSR_1/CLK MUX2X1_88/Y gnd vdd DFFPOSX1
XDFFPOSX1_58 INVX1_30/A DFFSR_8/CLK MUX2X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_69 INVX1_75/A CLKBUF1_3/Y MUX2X1_54/Y gnd vdd DFFPOSX1
XFILL_11_2_1 gnd vdd FILL
XNOR3X1_14 NOR3X1_14/A NOR3X1_14/B OAI22X1_6/Y gnd NOR3X1_14/Y vdd NOR3X1
XBUFX2_7 BUFX2_7/A gnd dout[6] vdd BUFX2
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XNAND2X1_2 INVX4_1/Y INVX1_43/A gnd MUX2X1_1/S vdd NAND2X1
XAOI21X1_7 NOR3X1_16/Y AOI21X1_7/B AOI21X1_7/C gnd DFFSR_7/D vdd AOI21X1
XFILL_8_2_1 gnd vdd FILL
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XFILL_0_1_1 gnd vdd FILL
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A OR2X2_2/Y gnd NOR2X1_5/Y vdd NOR2X1
XDFFPOSX1_2 INVX1_12/A CLKBUF1_3/Y MUX2X1_11/Y gnd vdd DFFPOSX1
XAOI21X1_26 INVX8_3/Y AND2X2_2/Y NOR2X1_39/Y gnd AOI21X1_26/Y vdd AOI21X1
XAOI21X1_15 INVX8_8/Y AND2X2_1/Y NOR2X1_26/Y gnd AOI21X1_15/Y vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XDFFPOSX1_15 INVX1_9/A CLKBUF1_8/Y MUX2X1_8/Y gnd vdd DFFPOSX1
XDFFPOSX1_59 INVX1_34/A DFFSR_1/CLK MUX2X1_60/Y gnd vdd DFFPOSX1
XDFFPOSX1_37 INVX1_99/A CLKBUF1_7/Y MUX2X1_84/Y gnd vdd DFFPOSX1
XDFFPOSX1_48 INVX1_94/A CLKBUF1_3/Y MUX2X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 INVX1_28/A DFFSR_8/CLK MUX2X1_89/Y gnd vdd DFFPOSX1
XNOR3X1_15 NOR3X1_15/A NOR3X1_15/B NOR3X1_15/C gnd AOI21X1_6/B vdd NOR3X1
XBUFX2_8 BUFX2_8/A gnd dout[7] vdd BUFX2
XNAND2X1_3 addr[0] INVX1_2/Y gnd INVX4_3/A vdd NAND2X1
XAOI21X1_8 NOR3X1_18/Y NOR3X1_19/Y AOI21X1_8/C gnd DFFSR_8/D vdd AOI21X1
XMUX2X1_100 INVX1_42/Y INVX8_6/Y MUX2X1_1/S gnd MUX2X1_100/Y vdd MUX2X1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XDFFPOSX1_3 INVX1_13/A CLKBUF1_2/Y MUX2X1_12/Y gnd vdd DFFPOSX1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XNOR2X1_6 OR2X2_2/Y INVX2_3/A gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_27 INVX8_4/Y AND2X2_2/Y NOR2X1_40/Y gnd AOI21X1_27/Y vdd AOI21X1
XAOI21X1_16 INVX8_1/Y AND2X2_1/Y NOR2X1_27/Y gnd AOI21X1_16/Y vdd AOI21X1
XDFFPOSX1_27 INVX1_32/A CLKBUF1_4/Y MUX2X1_90/Y gnd vdd DFFPOSX1
XDFFPOSX1_16 INVX1_10/A CLKBUF1_3/Y MUX2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 INVX1_100/A CLKBUF1_5/Y MUX2X1_85/Y gnd vdd DFFPOSX1
XDFFPOSX1_49 INVX1_79/A CLKBUF1_1/Y MUX2X1_64/Y gnd vdd DFFPOSX1
XFILL_14_2_0 gnd vdd FILL
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XNOR3X1_16 NOR3X1_16/A NOR3X1_16/B NOR3X1_16/C gnd NOR3X1_16/Y vdd NOR3X1
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XAOI21X1_9 INVX8_2/Y AND2X2_1/Y AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XNAND2X1_4 INVX4_1/Y NOR2X1_1/Y gnd MUX2X1_10/S vdd NAND2X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XMUX2X1_101 INVX1_109/Y INVX8_7/Y MUX2X1_1/S gnd MUX2X1_101/Y vdd MUX2X1
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XDFFPOSX1_4 INVX1_14/A CLKBUF1_10/Y MUX2X1_13/Y gnd vdd DFFPOSX1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XNOR2X1_7 INVX4_3/A INVX2_2/A gnd NOR2X1_7/Y vdd NOR2X1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XAOI21X1_28 INVX8_5/Y AND2X2_2/Y NOR2X1_41/Y gnd AOI21X1_28/Y vdd AOI21X1
XAOI21X1_17 INVX8_2/Y MUX2X1_18/S NOR2X1_29/Y gnd AOI21X1_17/Y vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XDFFPOSX1_28 INVX1_36/A DFFSR_1/CLK MUX2X1_91/Y gnd vdd DFFPOSX1
XDFFPOSX1_39 INVX1_101/A CLKBUF1_5/Y MUX2X1_86/Y gnd vdd DFFPOSX1
XDFFPOSX1_17 INVX1_105/A CLKBUF1_9/Y MUX2X1_96/Y gnd vdd DFFPOSX1
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd MUX2X1_85/A vdd INVX1
XNOR3X1_17 NOR3X1_17/A NOR3X1_17/B NOR3X1_17/C gnd AOI21X1_7/B vdd NOR3X1
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XMUX2X1_90 INVX1_32/Y INVX8_4/Y MUX2X1_91/S gnd MUX2X1_90/Y vdd MUX2X1
XNAND2X1_5 addr[0] addr[1] gnd INVX2_1/A vdd NAND2X1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XDFFPOSX1_5 INVX1_15/A CLKBUF1_3/Y MUX2X1_14/Y gnd vdd DFFPOSX1
XMUX2X1_102 INVX1_110/Y INVX8_8/Y MUX2X1_1/S gnd MUX2X1_102/Y vdd MUX2X1
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XAOI21X1_29 INVX8_6/Y AND2X2_2/Y NOR2X1_42/Y gnd AOI21X1_29/Y vdd AOI21X1
XNOR2X1_8 NOR2X1_8/A INVX2_2/A gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_18 INVX8_3/Y MUX2X1_18/S NOR2X1_30/Y gnd AOI21X1_18/Y vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XDFFPOSX1_29 INVX1_103/A CLKBUF1_3/Y MUX2X1_92/Y gnd vdd DFFPOSX1
XDFFPOSX1_18 INVX1_106/A CLKBUF1_7/Y MUX2X1_97/Y gnd vdd DFFPOSX1
XINVX1_101 INVX1_101/A gnd INVX1_101/Y vdd INVX1
XNOR3X1_18 NOR3X1_18/A NOR3X1_18/B NOR3X1_18/C gnd NOR3X1_18/Y vdd NOR3X1
XNOR2X1_40 NOR2X1_40/A AND2X2_2/Y gnd NOR2X1_40/Y vdd NOR2X1
XNAND2X1_6 addr[2] NOR3X1_4/A gnd INVX2_2/A vdd NAND2X1
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XMUX2X1_80 INVX1_95/Y INVX8_2/Y MUX2X1_80/S gnd MUX2X1_80/Y vdd MUX2X1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XMUX2X1_91 INVX1_36/Y INVX8_5/Y MUX2X1_91/S gnd MUX2X1_91/Y vdd MUX2X1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XDFFPOSX1_6 INVX1_16/A CLKBUF1_3/Y MUX2X1_15/Y gnd vdd DFFPOSX1
XNOR2X1_9 OR2X2_2/Y INVX2_2/A gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 INVX8_4/Y MUX2X1_18/S NOR2X1_31/Y gnd AOI21X1_19/Y vdd AOI21X1
XFILL_8_1 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XDFFPOSX1_19 AOI22X1_7/B CLKBUF1_9/Y MUX2X1_98/Y gnd vdd DFFPOSX1
XINVX1_102 INVX1_102/A gnd INVX1_102/Y vdd INVX1
XFILL_14_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XNOR3X1_19 NOR3X1_19/A NOR3X1_19/B NOR3X1_19/C gnd NOR3X1_19/Y vdd NOR3X1
XNOR2X1_41 NOR2X1_41/A AND2X2_2/Y gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_30 NOR2X1_30/A MUX2X1_18/S gnd NOR2X1_30/Y vdd NOR2X1
XNAND3X1_30 NAND2X1_52/Y NAND3X1_30/B NAND3X1_30/C gnd NOR3X1_19/B vdd NAND3X1
XNAND2X1_7 INVX2_1/Y INVX2_2/Y gnd OAI22X1_4/C vdd NAND2X1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XMUX2X1_70 INVX1_85/Y INVX8_8/Y MUX2X1_70/S gnd MUX2X1_70/Y vdd MUX2X1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XMUX2X1_92 MUX2X1_92/A INVX8_6/Y MUX2X1_91/S gnd MUX2X1_92/Y vdd MUX2X1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XMUX2X1_81 INVX1_96/Y INVX8_3/Y MUX2X1_80/S gnd MUX2X1_81/Y vdd MUX2X1
XDFFPOSX1_7 INVX1_17/A CLKBUF1_10/Y MUX2X1_16/Y gnd vdd DFFPOSX1
XFILL_1_2_1 gnd vdd FILL
XINVX1_103 INVX1_103/A gnd MUX2X1_92/A vdd INVX1
XFILL_14_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_20 NOR2X1_20/A AND2X2_1/Y gnd AOI21X1_9/C vdd NOR2X1
XNOR2X1_42 NOR2X1_42/A AND2X2_2/Y gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_31 NOR2X1_31/A MUX2X1_18/S gnd NOR2X1_31/Y vdd NOR2X1
XNAND3X1_31 NAND2X1_53/Y NAND3X1_31/B NAND3X1_31/C gnd NOR3X1_19/A vdd NAND3X1
XNAND3X1_20 NAND3X1_20/A NAND2X1_38/Y NAND2X1_39/Y gnd NOR3X1_13/A vdd NAND3X1
XMUX2X1_60 INVX8_4/Y INVX1_34/Y NOR2X1_48/B gnd MUX2X1_60/Y vdd MUX2X1
XMUX2X1_82 INVX1_97/Y INVX8_4/Y MUX2X1_80/S gnd MUX2X1_82/Y vdd MUX2X1
XNAND2X1_8 addr[3] addr[2] gnd NOR2X1_5/A vdd NAND2X1
XMUX2X1_71 INVX1_86/Y INVX8_1/Y MUX2X1_70/S gnd MUX2X1_71/Y vdd MUX2X1
XMUX2X1_93 INVX1_46/Y INVX8_7/Y MUX2X1_91/S gnd MUX2X1_93/Y vdd MUX2X1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XDFFPOSX1_8 INVX1_18/A CLKBUF1_10/Y MUX2X1_17/Y gnd vdd DFFPOSX1
XINVX1_23 addr[3] gnd NOR3X1_4/A vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_104 INVX1_104/A gnd MUX2X1_95/A vdd INVX1
XNOR2X1_43 NOR2X1_43/A AND2X2_2/Y gnd NOR2X1_43/Y vdd NOR2X1
XNAND3X1_10 NAND3X1_9/Y NAND2X1_24/Y NAND3X1_10/C gnd NOR3X1_9/A vdd NAND3X1
XNAND3X1_21 INVX1_8/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_21/Y vdd NAND3X1
XNOR2X1_32 NOR2X1_32/A MUX2X1_18/S gnd NOR2X1_32/Y vdd NOR2X1
XNOR2X1_10 INVX4_3/A INVX2_3/A gnd INVX1_45/A vdd NOR2X1
XNOR2X1_21 AOI22X1_6/A AND2X2_1/Y gnd NOR2X1_21/Y vdd NOR2X1
XMUX2X1_83 INVX1_98/Y INVX8_5/Y MUX2X1_80/S gnd MUX2X1_83/Y vdd MUX2X1
XMUX2X1_61 INVX8_5/Y INVX1_38/Y NOR2X1_48/B gnd MUX2X1_61/Y vdd MUX2X1
XMUX2X1_50 INVX1_71/Y INVX8_2/Y MUX2X1_52/S gnd MUX2X1_50/Y vdd MUX2X1
XMUX2X1_72 INVX1_87/Y INVX8_2/Y MUX2X1_77/S gnd MUX2X1_72/Y vdd MUX2X1
XNAND2X1_9 addr[1] NOR3X1_2/A gnd NOR2X1_8/A vdd NAND2X1
XMUX2X1_94 INVX1_50/Y INVX8_8/Y MUX2X1_91/S gnd MUX2X1_94/Y vdd MUX2X1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XDFFPOSX1_9 INVX1_3/A CLKBUF1_8/Y MUX2X1_2/Y gnd vdd DFFPOSX1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 addr[0] gnd NOR3X1_2/A vdd INVX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XFILL_12_1_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XFILL_6_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XINVX1_105 INVX1_105/A gnd MUX2X1_96/A vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XNOR2X1_44 NOR2X1_44/A AND2X2_2/Y gnd NOR2X1_44/Y vdd NOR2X1
XNAND3X1_22 NAND3X1_21/Y NAND3X1_22/B NAND3X1_22/C gnd NOR3X1_15/A vdd NAND3X1
XNAND3X1_11 NAND3X1_11/A NAND2X1_28/Y AOI22X1_9/Y gnd NOR3X1_9/B vdd NAND3X1
XNOR2X1_22 AOI22X1_9/A AND2X2_1/Y gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_11 INVX2_1/A NOR2X1_5/A gnd AND2X2_1/A vdd NOR2X1
XNOR2X1_33 NOR2X1_33/A MUX2X1_18/S gnd NOR2X1_33/Y vdd NOR2X1
XMUX2X1_73 INVX1_88/Y INVX8_3/Y MUX2X1_77/S gnd MUX2X1_73/Y vdd MUX2X1
XMUX2X1_84 INVX1_99/Y INVX8_6/Y MUX2X1_80/S gnd MUX2X1_84/Y vdd MUX2X1
XMUX2X1_40 INVX1_53/Y INVX8_8/Y OR2X2_3/Y gnd MUX2X1_40/Y vdd MUX2X1
XMUX2X1_95 MUX2X1_95/A INVX8_1/Y MUX2X1_91/S gnd MUX2X1_95/Y vdd MUX2X1
XMUX2X1_51 INVX1_72/Y INVX8_3/Y MUX2X1_52/S gnd MUX2X1_51/Y vdd MUX2X1
XMUX2X1_62 INVX8_7/Y INVX1_48/Y NOR2X1_48/B gnd MUX2X1_62/Y vdd MUX2X1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XFILL_12_1_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XCLKBUF1_10 clk gnd CLKBUF1_10/Y vdd CLKBUF1
XFILL_1_0_1 gnd vdd FILL
XFILL_9_1_1 gnd vdd FILL
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XNAND3X1_12 INVX1_6/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_13/B vdd NAND3X1
XNAND3X1_23 NAND3X1_23/A NAND2X1_45/Y AOI22X1_17/Y gnd NOR3X1_15/B vdd NAND3X1
XNOR2X1_12 NOR2X1_5/A NOR2X1_8/A gnd INVX2_5/A vdd NOR2X1
XMUX2X1_52 INVX1_73/Y INVX8_4/Y MUX2X1_52/S gnd MUX2X1_52/Y vdd MUX2X1
XMUX2X1_30 INVX1_61/Y INVX8_6/Y MUX2X1_29/S gnd MUX2X1_30/Y vdd MUX2X1
XMUX2X1_41 INVX1_55/Y INVX8_1/Y OR2X2_3/Y gnd MUX2X1_41/Y vdd MUX2X1
XNOR2X1_34 NOR2X1_34/A MUX2X1_18/S gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A AND2X2_1/Y gnd NOR2X1_23/Y vdd NOR2X1
XMUX2X1_63 INVX8_8/Y INVX1_52/Y NOR2X1_48/B gnd MUX2X1_63/Y vdd MUX2X1
XNOR2X1_45 NOR2X1_45/A AND2X2_2/Y gnd NOR2X1_45/Y vdd NOR2X1
XMUX2X1_74 INVX1_89/Y INVX8_4/Y MUX2X1_77/S gnd MUX2X1_74/Y vdd MUX2X1
XMUX2X1_85 MUX2X1_85/A INVX8_7/Y MUX2X1_80/S gnd MUX2X1_85/Y vdd MUX2X1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XINVX1_26 NOR2X1_8/A gnd INVX1_26/Y vdd INVX1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XMUX2X1_96 MUX2X1_96/A INVX8_2/Y MUX2X1_1/S gnd MUX2X1_96/Y vdd MUX2X1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XOAI21X1_10 INVX1_45/Y INVX1_44/Y NAND2X1_34/Y gnd NOR3X1_12/A vdd OAI21X1
XCLKBUF1_11 clk gnd DFFSR_1/CLK vdd CLKBUF1
XINVX1_107 AOI22X1_7/B gnd MUX2X1_98/A vdd INVX1
XFILL_10_2_0 gnd vdd FILL
XNAND3X1_13 NAND2X1_30/Y NAND3X1_13/B NAND3X1_13/C gnd NOR3X1_11/A vdd NAND3X1
XNAND3X1_24 INVX1_9/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_24/Y vdd NAND3X1
XNOR2X1_13 BUFX2_2/A NOR2X1_3/B gnd AOI21X1_2/C vdd NOR2X1
XNOR2X1_24 NOR2X1_24/A AND2X2_1/Y gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_46 INVX4_1/A OAI22X1_4/C gnd NOR2X1_48/B vdd NOR2X1
XNOR2X1_35 INVX4_1/A INVX4_5/Y gnd MUX2X1_20/S vdd NOR2X1
XFILL_16_1 gnd vdd FILL
XDFFSR_1 DFFSR_1/Q DFFSR_1/CLK rst_n vdd DFFSR_1/D gnd vdd DFFSR
XMUX2X1_75 INVX1_90/Y INVX8_5/Y MUX2X1_77/S gnd MUX2X1_75/Y vdd MUX2X1
XMUX2X1_42 INVX1_65/Y INVX8_2/Y MUX2X1_45/S gnd MUX2X1_42/Y vdd MUX2X1
XMUX2X1_20 INVX8_2/Y INVX1_21/Y MUX2X1_20/S gnd MUX2X1_20/Y vdd MUX2X1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XMUX2X1_86 INVX1_101/Y INVX8_8/Y MUX2X1_80/S gnd MUX2X1_86/Y vdd MUX2X1
XMUX2X1_31 INVX1_62/Y INVX8_7/Y MUX2X1_29/S gnd MUX2X1_31/Y vdd MUX2X1
XMUX2X1_53 INVX1_74/Y INVX8_5/Y MUX2X1_52/S gnd MUX2X1_53/Y vdd MUX2X1
XINVX1_27 addr[2] gnd INVX1_27/Y vdd INVX1
XMUX2X1_64 INVX1_79/Y INVX8_2/Y MUX2X1_70/S gnd MUX2X1_64/Y vdd MUX2X1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XMUX2X1_97 INVX1_106/Y INVX8_3/Y MUX2X1_1/S gnd MUX2X1_97/Y vdd MUX2X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_11 INVX4_4/Y INVX1_46/Y NOR2X1_3/B gnd NOR3X1_14/B vdd OAI21X1
XFILL_4_0_0 gnd vdd FILL
XINVX1_108 INVX1_108/A gnd MUX2X1_99/A vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNOR2X1_14 DFFSR_3/Q NOR2X1_3/B gnd AOI21X1_3/C vdd NOR2X1
XNAND3X1_25 NAND3X1_25/A NAND3X1_24/Y NAND3X1_25/C gnd NOR3X1_17/A vdd NAND3X1
XNOR2X1_36 NOR2X1_36/A MUX2X1_20/S gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_14 INVX1_74/A INVX2_4/Y INVX2_3/Y gnd NAND3X1_14/Y vdd NAND3X1
XNOR2X1_47 NOR2X1_47/A NOR2X1_48/B gnd NOR2X1_47/Y vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A AND2X2_1/Y gnd NOR2X1_25/Y vdd NOR2X1
XDFFSR_2 BUFX2_2/A DFFSR_1/CLK rst_n vdd DFFSR_2/D gnd vdd DFFSR
XMUX2X1_10 INVX1_11/Y INVX8_2/Y MUX2X1_10/S gnd MUX2X1_10/Y vdd MUX2X1
XMUX2X1_21 INVX8_3/Y INVX1_29/Y MUX2X1_20/S gnd MUX2X1_21/Y vdd MUX2X1
XMUX2X1_32 INVX1_63/Y INVX8_8/Y MUX2X1_29/S gnd MUX2X1_32/Y vdd MUX2X1
XMUX2X1_65 INVX1_80/Y INVX8_3/Y MUX2X1_70/S gnd MUX2X1_65/Y vdd MUX2X1
XMUX2X1_98 MUX2X1_98/A INVX8_4/Y MUX2X1_1/S gnd MUX2X1_98/Y vdd MUX2X1
XMUX2X1_76 INVX1_91/Y INVX8_6/Y MUX2X1_77/S gnd MUX2X1_76/Y vdd MUX2X1
XMUX2X1_43 INVX1_66/Y INVX8_3/Y MUX2X1_45/S gnd MUX2X1_43/Y vdd MUX2X1
XMUX2X1_54 INVX1_75/Y INVX8_6/Y MUX2X1_52/S gnd MUX2X1_54/Y vdd MUX2X1
XMUX2X1_87 INVX1_102/Y INVX8_1/Y MUX2X1_80/S gnd MUX2X1_87/Y vdd MUX2X1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_12 OR2X2_3/A INVX1_49/Y NAND2X1_40/Y gnd NOR3X1_14/A vdd OAI21X1
XFILL_4_0_1 gnd vdd FILL
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XNOR2X1_15 BUFX2_4/A NOR2X1_3/B gnd AOI21X1_4/C vdd NOR2X1
XNOR2X1_26 NOR2X1_26/A AND2X2_1/Y gnd NOR2X1_26/Y vdd NOR2X1
XNAND3X1_15 NAND3X1_14/Y NAND3X1_15/B AOI22X1_12/Y gnd NOR3X1_11/B vdd NAND3X1
XNAND3X1_26 INVX1_77/A INVX2_4/Y INVX2_3/Y gnd NAND3X1_27/A vdd NAND3X1
XNOR2X1_37 NOR2X1_37/A MUX2X1_20/S gnd NOR2X1_37/Y vdd NOR2X1
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XDFFSR_3 DFFSR_3/Q DFFSR_1/CLK rst_n vdd DFFSR_3/D gnd vdd DFFSR
XMUX2X1_77 INVX1_92/Y INVX8_7/Y MUX2X1_77/S gnd MUX2X1_77/Y vdd MUX2X1
XMUX2X1_88 INVX1_20/Y INVX8_2/Y MUX2X1_91/S gnd MUX2X1_88/Y vdd MUX2X1
XMUX2X1_44 INVX1_67/Y INVX8_4/Y MUX2X1_45/S gnd MUX2X1_44/Y vdd MUX2X1
XMUX2X1_55 INVX1_76/Y INVX8_7/Y MUX2X1_52/S gnd MUX2X1_55/Y vdd MUX2X1
XMUX2X1_22 INVX8_4/Y INVX1_33/Y MUX2X1_20/S gnd MUX2X1_22/Y vdd MUX2X1
XMUX2X1_33 INVX1_64/Y INVX8_1/Y MUX2X1_29/S gnd MUX2X1_33/Y vdd MUX2X1
XMUX2X1_66 INVX1_81/Y INVX8_4/Y MUX2X1_70/S gnd MUX2X1_66/Y vdd MUX2X1
XMUX2X1_99 MUX2X1_99/A INVX8_5/Y MUX2X1_1/S gnd MUX2X1_99/Y vdd MUX2X1
XMUX2X1_11 INVX1_12/Y INVX8_3/Y MUX2X1_10/S gnd MUX2X1_11/Y vdd MUX2X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XOAI21X1_13 INVX4_4/Y INVX1_50/Y NOR2X1_3/B gnd NOR3X1_16/B vdd OAI21X1
XFILL_13_2_0 gnd vdd FILL
XNOR2X1_38 NOR2X1_38/A AND2X2_2/Y gnd NOR2X1_38/Y vdd NOR2X1
XNOR2X1_16 BUFX2_5/A NOR2X1_3/B gnd AOI21X1_5/C vdd NOR2X1
XNOR2X1_27 NOR2X1_27/A AND2X2_1/Y gnd NOR2X1_27/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNAND3X1_27 NAND3X1_27/A NAND2X1_50/Y AOI22X1_20/Y gnd NOR3X1_17/B vdd NAND3X1
XNAND3X1_16 NOR2X1_47/A INVX2_1/Y INVX2_2/Y gnd NAND3X1_18/A vdd NAND3X1
XMUX2X1_45 INVX1_68/Y INVX8_5/Y MUX2X1_45/S gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_78 INVX1_93/Y INVX8_8/Y MUX2X1_77/S gnd MUX2X1_78/Y vdd MUX2X1
XMUX2X1_34 INVX1_25/Y INVX8_2/Y OR2X2_3/Y gnd MUX2X1_34/Y vdd MUX2X1
XMUX2X1_23 INVX8_5/Y INVX1_37/Y MUX2X1_20/S gnd MUX2X1_23/Y vdd MUX2X1
XMUX2X1_12 INVX1_13/Y INVX8_4/Y MUX2X1_10/S gnd MUX2X1_12/Y vdd MUX2X1
XFILL_10_0_0 gnd vdd FILL
XMUX2X1_67 INVX1_82/Y INVX8_5/Y MUX2X1_70/S gnd MUX2X1_67/Y vdd MUX2X1
XMUX2X1_56 INVX1_77/Y INVX8_8/Y MUX2X1_52/S gnd MUX2X1_56/Y vdd MUX2X1
XMUX2X1_89 INVX1_28/Y INVX8_3/Y MUX2X1_91/S gnd MUX2X1_89/Y vdd MUX2X1
XDFFSR_4 BUFX2_4/A DFFSR_1/CLK rst_n vdd DFFSR_4/D gnd vdd DFFSR
XINVX1_19 re gnd NOR2X1_2/B vdd INVX1
XNAND2X1_60 INVX4_1/Y NOR2X1_7/Y gnd MUX2X1_77/S vdd NAND2X1
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_14 OR2X2_3/A INVX1_53/Y NAND2X1_46/Y gnd NOR3X1_16/A vdd OAI21X1
XDFFPOSX1_120 INVX1_54/A CLKBUF1_1/Y MUX2X1_19/Y gnd vdd DFFPOSX1
XFILL_13_2_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_2_1 gnd vdd FILL
XAND2X2_1 AND2X2_1/A INVX4_1/Y gnd AND2X2_1/Y vdd AND2X2
XNAND3X1_17 INVX1_7/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_18/B vdd NAND3X1
XNOR2X1_17 BUFX2_6/A NOR2X1_3/B gnd AOI21X1_6/C vdd NOR2X1
XNOR2X1_28 INVX4_1/A INVX2_5/Y gnd MUX2X1_18/S vdd NOR2X1
XNAND3X1_28 NOR2X1_48/A INVX2_1/Y INVX2_2/Y gnd NAND3X1_30/B vdd NAND3X1
XNOR2X1_39 NOR2X1_39/A AND2X2_2/Y gnd NOR2X1_39/Y vdd NOR2X1
XFILL_10_0_1 gnd vdd FILL
XMUX2X1_57 INVX1_78/Y INVX8_1/Y MUX2X1_52/S gnd MUX2X1_57/Y vdd MUX2X1
XMUX2X1_35 INVX1_31/Y INVX8_3/Y OR2X2_3/Y gnd MUX2X1_35/Y vdd MUX2X1
XMUX2X1_68 INVX1_83/Y INVX8_6/Y MUX2X1_70/S gnd MUX2X1_68/Y vdd MUX2X1
XMUX2X1_13 INVX1_14/Y INVX8_5/Y MUX2X1_10/S gnd MUX2X1_13/Y vdd MUX2X1
XFILL_2_1_1 gnd vdd FILL
XMUX2X1_46 INVX1_44/Y INVX8_6/Y MUX2X1_45/S gnd MUX2X1_46/Y vdd MUX2X1
XMUX2X1_79 INVX1_94/Y INVX8_1/Y MUX2X1_77/S gnd MUX2X1_79/Y vdd MUX2X1
XMUX2X1_24 INVX8_7/Y INVX1_47/Y MUX2X1_20/S gnd MUX2X1_24/Y vdd MUX2X1
XDFFSR_5 BUFX2_5/A CLKBUF1_4/Y rst_n vdd DFFSR_5/D gnd vdd DFFSR
XNAND2X1_50 NOR2X1_34/A INVX2_5/A gnd NAND2X1_50/Y vdd NAND2X1
XNAND2X1_61 INVX4_1/Y NOR2X1_9/Y gnd MUX2X1_80/S vdd NAND2X1
XOAI21X1_15 INVX2_5/Y INVX1_54/Y NOR2X1_3/B gnd NOR3X1_18/B vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XDFFPOSX1_121 NOR2X1_20/A CLKBUF1_2/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_110 INVX1_47/A DFFSR_8/CLK MUX2X1_24/Y gnd vdd DFFPOSX1
XINVX1_2 addr[1] gnd INVX1_2/Y vdd INVX1
XAND2X2_2 AND2X2_2/A INVX4_1/Y gnd AND2X2_2/Y vdd AND2X2
XNAND3X1_29 INVX1_10/A INVX4_2/Y INVX4_3/Y gnd NAND3X1_30/C vdd NAND3X1
XNOR2X1_18 BUFX2_7/A NOR2X1_3/B gnd AOI21X1_7/C vdd NOR2X1
XNAND3X1_18 NAND3X1_18/A NAND3X1_18/B NAND2X1_35/Y gnd NOR3X1_13/B vdd NAND3X1
XNOR2X1_29 NOR2X1_29/A MUX2X1_18/S gnd NOR2X1_29/Y vdd NOR2X1
XMUX2X1_36 INVX1_35/Y INVX8_4/Y OR2X2_3/Y gnd MUX2X1_36/Y vdd MUX2X1
XMUX2X1_47 INVX1_69/Y INVX8_7/Y MUX2X1_45/S gnd MUX2X1_47/Y vdd MUX2X1
XMUX2X1_58 INVX8_2/Y INVX1_22/Y NOR2X1_48/B gnd MUX2X1_58/Y vdd MUX2X1
XDFFSR_6 BUFX2_6/A CLKBUF1_4/Y rst_n vdd DFFSR_6/D gnd vdd DFFSR
XMUX2X1_69 INVX1_84/Y INVX8_7/Y MUX2X1_70/S gnd MUX2X1_69/Y vdd MUX2X1
XNAND2X1_40 INVX1_62/A NOR2X1_5/Y gnd NAND2X1_40/Y vdd NAND2X1
XNAND2X1_51 INVX1_86/A NOR2X1_8/Y gnd NAND2X1_51/Y vdd NAND2X1
XMUX2X1_14 INVX1_15/Y INVX8_6/Y MUX2X1_10/S gnd MUX2X1_14/Y vdd MUX2X1
XNAND2X1_62 INVX4_1/Y INVX4_4/A gnd MUX2X1_91/S vdd NAND2X1
XMUX2X1_25 INVX8_8/Y INVX1_51/Y MUX2X1_20/S gnd MUX2X1_25/Y vdd MUX2X1
XOAI21X1_16 INVX1_45/Y INVX1_56/Y NAND2X1_51/Y gnd NOR3X1_18/A vdd OAI21X1
XDFFPOSX1_100 INVX1_60/A CLKBUF1_4/Y MUX2X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 AOI22X1_6/A CLKBUF1_3/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_111 INVX1_51/A DFFSR_8/CLK MUX2X1_25/Y gnd vdd DFFPOSX1
XFILL_0_2_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XOR2X2_1 addr[3] addr[2] gnd INVX4_2/A vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_13_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XNAND3X1_19 NAND2X1_36/Y NAND3X1_19/B NAND3X1_19/C gnd NOR3X1_13/C vdd NAND3X1
XNOR2X1_19 BUFX2_8/A NOR2X1_3/B gnd AOI21X1_8/C vdd NOR2X1
XMUX2X1_48 INVX1_70/Y INVX8_8/Y MUX2X1_45/S gnd MUX2X1_48/Y vdd MUX2X1
XMUX2X1_37 INVX1_39/Y INVX8_5/Y OR2X2_3/Y gnd MUX2X1_37/Y vdd MUX2X1
XDFFSR_7 BUFX2_7/A CLKBUF1_4/Y rst_n vdd DFFSR_7/D gnd vdd DFFSR
XMUX2X1_26 INVX1_57/Y INVX8_2/Y MUX2X1_29/S gnd MUX2X1_26/Y vdd MUX2X1
XMUX2X1_59 INVX8_3/Y INVX1_30/Y NOR2X1_48/B gnd MUX2X1_59/Y vdd MUX2X1
XMUX2X1_15 INVX1_16/Y INVX8_7/Y MUX2X1_10/S gnd MUX2X1_15/Y vdd MUX2X1
XNAND2X1_30 NOR2X1_41/A AND2X2_2/A gnd NAND2X1_30/Y vdd NAND2X1
XNAND2X1_41 INVX1_76/A NOR2X1_6/Y gnd NAND3X1_22/B vdd NAND2X1
XNAND2X1_52 NOR2X1_45/A AND2X2_2/A gnd NAND2X1_52/Y vdd NAND2X1
XOAI22X1_1 INVX1_21/Y INVX4_5/Y OAI22X1_4/C INVX1_22/Y gnd NOR3X1_3/C vdd OAI22X1
XFILL_12_1 gnd vdd FILL
XDFFPOSX1_101 INVX1_61/A CLKBUF1_4/Y MUX2X1_30/Y gnd vdd DFFPOSX1
XDFFPOSX1_123 AOI22X1_9/A CLKBUF1_7/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XFILL_0_2_1 gnd vdd FILL
XDFFPOSX1_112 NOR2X1_37/A CLKBUF1_1/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XFILL_16_2_1 gnd vdd FILL
XOR2X2_2 addr[0] addr[1] gnd OR2X2_2/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XMUX2X1_27 INVX1_58/Y INVX8_3/Y MUX2X1_29/S gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_16 INVX1_17/Y INVX8_8/Y MUX2X1_10/S gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_49 INVX1_56/Y INVX8_1/Y MUX2X1_45/S gnd MUX2X1_49/Y vdd MUX2X1
XMUX2X1_38 INVX1_41/Y INVX8_6/Y OR2X2_3/Y gnd MUX2X1_38/Y vdd MUX2X1
XDFFSR_8 BUFX2_8/A DFFSR_8/CLK rst_n vdd DFFSR_8/D gnd vdd DFFSR
XNAND2X1_31 INVX1_90/A NOR2X1_7/Y gnd NAND3X1_13/C vdd NAND2X1
XNAND2X1_20 INVX1_88/A NOR2X1_7/Y gnd NAND3X1_6/C vdd NAND2X1
XNAND2X1_42 INVX1_92/A NOR2X1_7/Y gnd NAND3X1_22/C vdd NAND2X1
XNAND2X1_53 INVX1_18/A NOR2X1_1/Y gnd NAND2X1_53/Y vdd NAND2X1
XOAI22X1_2 INVX1_29/Y INVX4_5/Y OAI22X1_4/C INVX1_30/Y gnd NOR3X1_6/C vdd OAI22X1
XDFFPOSX1_102 INVX1_62/A CLKBUF1_1/Y MUX2X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_124 NOR2X1_23/A CLKBUF1_10/Y AOI21X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 NOR2X1_29/A CLKBUF1_7/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOR2X2_3 OR2X2_3/A INVX4_1/A gnd OR2X2_3/Y vdd OR2X2
.ends

